// weights_and_biases.vh

//initial begin
task initialize_weights_and_biases;
    weight_rom[0][0] = -32'd1644;
    weight_rom[0][1] = -32'd6462;
    weight_rom[0][2] = 32'd5716;
    weight_rom[0][3] = 32'd3081;
    weight_rom[0][4] = 32'd5671;
    weight_rom[0][5] = -32'd6290;
    weight_rom[0][6] = -32'd2069;
    weight_rom[0][7] = -32'd2711;
    weight_rom[0][8] = 32'd5823;
    weight_rom[0][9] = 32'd2588;
    weight_rom[0][10] = 32'd1548;
    weight_rom[0][11] = 32'd1118;
    weight_rom[0][12] = -32'd4179;
    weight_rom[0][13] = 32'd6450;
    weight_rom[0][14] = 32'd160;
    weight_rom[0][15] = 32'd2564;
    weight_rom[0][16] = 32'd570;
    weight_rom[0][17] = -32'd2893;
    weight_rom[0][18] = 32'd5659;
    weight_rom[0][19] = 32'd6344;
    weight_rom[0][20] = 32'd3860;
    weight_rom[0][21] = -32'd93;
    weight_rom[0][22] = -32'd14;
    weight_rom[0][23] = 32'd3394;
    weight_rom[0][24] = -32'd2452;
    weight_rom[0][25] = 32'd699;
    weight_rom[0][26] = -32'd4714;
    weight_rom[0][27] = 32'd4;
    weight_rom[0][28] = -32'd1221;
    weight_rom[0][29] = 32'd2703;
    weight_rom[0][30] = 32'd413;
    weight_rom[0][31] = 32'd1158;
    weight_rom[0][32] = -32'd6374;
    weight_rom[0][33] = 32'd1089;
    weight_rom[0][34] = -32'd1125;
    weight_rom[0][35] = -32'd4437;
    weight_rom[0][36] = 32'd5980;
    weight_rom[0][37] = 32'd162;
    weight_rom[0][38] = -32'd2441;
    weight_rom[0][39] = -32'd2075;
    weight_rom[0][40] = -32'd2384;
    weight_rom[0][41] = -32'd565;
    weight_rom[0][42] = 32'd1002;
    weight_rom[0][43] = -32'd2487;
    weight_rom[0][44] = -32'd4107;
    weight_rom[0][45] = 32'd3435;
    weight_rom[0][46] = 32'd3942;
    weight_rom[0][47] = -32'd4817;
    weight_rom[0][48] = 32'd3711;
    weight_rom[0][49] = -32'd5693;
    weight_rom[0][50] = 32'd2414;
    weight_rom[0][51] = -32'd1764;
    weight_rom[0][52] = -32'd3261;
    weight_rom[0][53] = 32'd3004;
    weight_rom[0][54] = -32'd3924;
    weight_rom[0][55] = 32'd3722;
    weight_rom[0][56] = -32'd3114;
    weight_rom[0][57] = -32'd4475;
    weight_rom[0][58] = -32'd404;
    weight_rom[0][59] = 32'd2122;
    weight_rom[0][60] = 32'd5735;
    weight_rom[0][61] = -32'd3185;
    weight_rom[0][62] = 32'd127;
    weight_rom[0][63] = 32'd6103;
    weight_rom[1][0] = 32'd5907;
    weight_rom[1][1] = 32'd140;
    weight_rom[1][2] = 32'd2569;
    weight_rom[1][3] = 32'd3977;
    weight_rom[1][4] = 32'd4798;
    weight_rom[1][5] = -32'd2332;
    weight_rom[1][6] = 32'd4210;
    weight_rom[1][7] = 32'd5194;
    weight_rom[1][8] = -32'd337;
    weight_rom[1][9] = 32'd2361;
    weight_rom[1][10] = 32'd2653;
    weight_rom[1][11] = 32'd4826;
    weight_rom[1][12] = 32'd2373;
    weight_rom[1][13] = 32'd4606;
    weight_rom[1][14] = 32'd2362;
    weight_rom[1][15] = -32'd6511;
    weight_rom[1][16] = -32'd5482;
    weight_rom[1][17] = 32'd1872;
    weight_rom[1][18] = -32'd1349;
    weight_rom[1][19] = -32'd2773;
    weight_rom[1][20] = 32'd2714;
    weight_rom[1][21] = -32'd1254;
    weight_rom[1][22] = -32'd6394;
    weight_rom[1][23] = -32'd5209;
    weight_rom[1][24] = -32'd3000;
    weight_rom[1][25] = 32'd41;
    weight_rom[1][26] = 32'd2243;
    weight_rom[1][27] = 32'd2501;
    weight_rom[1][28] = -32'd2251;
    weight_rom[1][29] = 32'd1608;
    weight_rom[1][30] = -32'd6125;
    weight_rom[1][31] = -32'd1341;
    weight_rom[1][32] = -32'd5484;
    weight_rom[1][33] = 32'd3017;
    weight_rom[1][34] = 32'd6002;
    weight_rom[1][35] = -32'd370;
    weight_rom[1][36] = -32'd1616;
    weight_rom[1][37] = -32'd1981;
    weight_rom[1][38] = 32'd1777;
    weight_rom[1][39] = 32'd1945;
    weight_rom[1][40] = 32'd5565;
    weight_rom[1][41] = -32'd326;
    weight_rom[1][42] = -32'd2070;
    weight_rom[1][43] = -32'd4171;
    weight_rom[1][44] = -32'd4086;
    weight_rom[1][45] = 32'd5717;
    weight_rom[1][46] = -32'd640;
    weight_rom[1][47] = 32'd614;
    weight_rom[1][48] = -32'd4350;
    weight_rom[1][49] = 32'd647;
    weight_rom[1][50] = 32'd5012;
    weight_rom[1][51] = 32'd4477;
    weight_rom[1][52] = -32'd2351;
    weight_rom[1][53] = 32'd4911;
    weight_rom[1][54] = -32'd3730;
    weight_rom[1][55] = -32'd1378;
    weight_rom[1][56] = -32'd3384;
    weight_rom[1][57] = -32'd164;
    weight_rom[1][58] = -32'd1733;
    weight_rom[1][59] = -32'd460;
    weight_rom[1][60] = 32'd391;
    weight_rom[1][61] = -32'd6279;
    weight_rom[1][62] = 32'd1117;
    weight_rom[1][63] = -32'd6358;
    weight_rom[2][0] = 32'd3040;
    weight_rom[2][1] = -32'd1082;
    weight_rom[2][2] = 32'd918;
    weight_rom[2][3] = -32'd2856;
    weight_rom[2][4] = -32'd5960;
    weight_rom[2][5] = -32'd3782;
    weight_rom[2][6] = -32'd5103;
    weight_rom[2][7] = -32'd6383;
    weight_rom[2][8] = 32'd4745;
    weight_rom[2][9] = 32'd1554;
    weight_rom[2][10] = 32'd781;
    weight_rom[2][11] = -32'd3855;
    weight_rom[2][12] = -32'd4175;
    weight_rom[2][13] = -32'd3820;
    weight_rom[2][14] = -32'd6007;
    weight_rom[2][15] = 32'd1567;
    weight_rom[2][16] = -32'd546;
    weight_rom[2][17] = 32'd2544;
    weight_rom[2][18] = -32'd5412;
    weight_rom[2][19] = 32'd6044;
    weight_rom[2][20] = -32'd5895;
    weight_rom[2][21] = 32'd405;
    weight_rom[2][22] = -32'd6435;
    weight_rom[2][23] = 32'd181;
    weight_rom[2][24] = 32'd1280;
    weight_rom[2][25] = -32'd4012;
    weight_rom[2][26] = 32'd1579;
    weight_rom[2][27] = 32'd2583;
    weight_rom[2][28] = -32'd603;
    weight_rom[2][29] = 32'd6423;
    weight_rom[2][30] = -32'd319;
    weight_rom[2][31] = 32'd6210;
    weight_rom[2][32] = -32'd3164;
    weight_rom[2][33] = -32'd1771;
    weight_rom[2][34] = 32'd538;
    weight_rom[2][35] = 32'd700;
    weight_rom[2][36] = -32'd2107;
    weight_rom[2][37] = -32'd1640;
    weight_rom[2][38] = -32'd1887;
    weight_rom[2][39] = -32'd5656;
    weight_rom[2][40] = -32'd5816;
    weight_rom[2][41] = -32'd1493;
    weight_rom[2][42] = 32'd4062;
    weight_rom[2][43] = 32'd54;
    weight_rom[2][44] = -32'd4138;
    weight_rom[2][45] = 32'd5776;
    weight_rom[2][46] = 32'd2866;
    weight_rom[2][47] = 32'd606;
    weight_rom[2][48] = 32'd160;
    weight_rom[2][49] = 32'd1190;
    weight_rom[2][50] = -32'd3886;
    weight_rom[2][51] = 32'd715;
    weight_rom[2][52] = -32'd4784;
    weight_rom[2][53] = 32'd5750;
    weight_rom[2][54] = -32'd2728;
    weight_rom[2][55] = 32'd1914;
    weight_rom[2][56] = -32'd222;
    weight_rom[2][57] = -32'd1781;
    weight_rom[2][58] = -32'd5234;
    weight_rom[2][59] = 32'd1711;
    weight_rom[2][60] = 32'd1506;
    weight_rom[2][61] = -32'd3629;
    weight_rom[2][62] = -32'd1843;
    weight_rom[2][63] = -32'd247;
    weight_rom[3][0] = 32'd1293;
    weight_rom[3][1] = -32'd3642;
    weight_rom[3][2] = -32'd5279;
    weight_rom[3][3] = -32'd4227;
    weight_rom[3][4] = -32'd6208;
    weight_rom[3][5] = -32'd2261;
    weight_rom[3][6] = 32'd4540;
    weight_rom[3][7] = -32'd5432;
    weight_rom[3][8] = 32'd4516;
    weight_rom[3][9] = 32'd3312;
    weight_rom[3][10] = -32'd6425;
    weight_rom[3][11] = -32'd5086;
    weight_rom[3][12] = 32'd329;
    weight_rom[3][13] = 32'd5643;
    weight_rom[3][14] = -32'd5442;
    weight_rom[3][15] = -32'd1894;
    weight_rom[3][16] = -32'd200;
    weight_rom[3][17] = 32'd165;
    weight_rom[3][18] = 32'd1534;
    weight_rom[3][19] = -32'd1448;
    weight_rom[3][20] = -32'd5598;
    weight_rom[3][21] = 32'd1246;
    weight_rom[3][22] = -32'd1873;
    weight_rom[3][23] = 32'd116;
    weight_rom[3][24] = 32'd4798;
    weight_rom[3][25] = 32'd4703;
    weight_rom[3][26] = 32'd3175;
    weight_rom[3][27] = 32'd1948;
    weight_rom[3][28] = 32'd3439;
    weight_rom[3][29] = -32'd2465;
    weight_rom[3][30] = -32'd1209;
    weight_rom[3][31] = 32'd579;
    weight_rom[3][32] = -32'd6188;
    weight_rom[3][33] = 32'd1847;
    weight_rom[3][34] = 32'd1377;
    weight_rom[3][35] = 32'd921;
    weight_rom[3][36] = -32'd5735;
    weight_rom[3][37] = 32'd1590;
    weight_rom[3][38] = -32'd4607;
    weight_rom[3][39] = 32'd5208;
    weight_rom[3][40] = -32'd188;
    weight_rom[3][41] = 32'd6117;
    weight_rom[3][42] = -32'd3430;
    weight_rom[3][43] = -32'd2322;
    weight_rom[3][44] = -32'd5806;
    weight_rom[3][45] = -32'd4262;
    weight_rom[3][46] = 32'd1130;
    weight_rom[3][47] = -32'd5380;
    weight_rom[3][48] = -32'd165;
    weight_rom[3][49] = 32'd2001;
    weight_rom[3][50] = 32'd4893;
    weight_rom[3][51] = 32'd5264;
    weight_rom[3][52] = -32'd2671;
    weight_rom[3][53] = 32'd3998;
    weight_rom[3][54] = -32'd4289;
    weight_rom[3][55] = -32'd4579;
    weight_rom[3][56] = 32'd5070;
    weight_rom[3][57] = 32'd1826;
    weight_rom[3][58] = -32'd2495;
    weight_rom[3][59] = -32'd660;
    weight_rom[3][60] = -32'd230;
    weight_rom[3][61] = -32'd5812;
    weight_rom[3][62] = -32'd322;
    weight_rom[3][63] = -32'd2184;
    weight_rom[4][0] = -32'd4508;
    weight_rom[4][1] = -32'd4982;
    weight_rom[4][2] = 32'd1507;
    weight_rom[4][3] = 32'd3284;
    weight_rom[4][4] = -32'd1619;
    weight_rom[4][5] = -32'd4983;
    weight_rom[4][6] = -32'd4882;
    weight_rom[4][7] = -32'd3828;
    weight_rom[4][8] = -32'd2371;
    weight_rom[4][9] = -32'd4474;
    weight_rom[4][10] = -32'd2274;
    weight_rom[4][11] = -32'd3017;
    weight_rom[4][12] = 32'd2739;
    weight_rom[4][13] = -32'd5028;
    weight_rom[4][14] = 32'd2835;
    weight_rom[4][15] = 32'd3856;
    weight_rom[4][16] = -32'd4380;
    weight_rom[4][17] = -32'd2551;
    weight_rom[4][18] = -32'd5061;
    weight_rom[4][19] = -32'd1500;
    weight_rom[4][20] = -32'd1273;
    weight_rom[4][21] = -32'd6423;
    weight_rom[4][22] = 32'd5586;
    weight_rom[4][23] = -32'd1713;
    weight_rom[4][24] = 32'd5855;
    weight_rom[4][25] = 32'd2319;
    weight_rom[4][26] = -32'd4326;
    weight_rom[4][27] = -32'd2945;
    weight_rom[4][28] = -32'd4902;
    weight_rom[4][29] = -32'd2097;
    weight_rom[4][30] = -32'd4440;
    weight_rom[4][31] = -32'd2945;
    weight_rom[4][32] = 32'd1721;
    weight_rom[4][33] = -32'd443;
    weight_rom[4][34] = -32'd3663;
    weight_rom[4][35] = -32'd3799;
    weight_rom[4][36] = -32'd181;
    weight_rom[4][37] = 32'd2866;
    weight_rom[4][38] = 32'd1264;
    weight_rom[4][39] = -32'd4988;
    weight_rom[4][40] = 32'd5410;
    weight_rom[4][41] = 32'd2584;
    weight_rom[4][42] = -32'd3612;
    weight_rom[4][43] = -32'd3170;
    weight_rom[4][44] = 32'd1150;
    weight_rom[4][45] = 32'd4911;
    weight_rom[4][46] = -32'd100;
    weight_rom[4][47] = -32'd1074;
    weight_rom[4][48] = 32'd1639;
    weight_rom[4][49] = -32'd3202;
    weight_rom[4][50] = -32'd5770;
    weight_rom[4][51] = 32'd5586;
    weight_rom[4][52] = 32'd947;
    weight_rom[4][53] = 32'd4595;
    weight_rom[4][54] = -32'd1581;
    weight_rom[4][55] = 32'd5670;
    weight_rom[4][56] = -32'd1594;
    weight_rom[4][57] = -32'd4862;
    weight_rom[4][58] = 32'd2146;
    weight_rom[4][59] = -32'd4081;
    weight_rom[4][60] = -32'd5326;
    weight_rom[4][61] = -32'd5198;
    weight_rom[4][62] = -32'd1788;
    weight_rom[4][63] = -32'd666;
    weight_rom[5][0] = -32'd4508;
    weight_rom[5][1] = -32'd2128;
    weight_rom[5][2] = 32'd6423;
    weight_rom[5][3] = 32'd4021;
    weight_rom[5][4] = 32'd4070;
    weight_rom[5][5] = 32'd5118;
    weight_rom[5][6] = -32'd1346;
    weight_rom[5][7] = -32'd6205;
    weight_rom[5][8] = 32'd4311;
    weight_rom[5][9] = 32'd4992;
    weight_rom[5][10] = 32'd232;
    weight_rom[5][11] = -32'd5805;
    weight_rom[5][12] = -32'd5152;
    weight_rom[5][13] = 32'd4160;
    weight_rom[5][14] = -32'd5608;
    weight_rom[5][15] = -32'd5334;
    weight_rom[5][16] = 32'd5841;
    weight_rom[5][17] = -32'd3766;
    weight_rom[5][18] = -32'd2028;
    weight_rom[5][19] = -32'd2092;
    weight_rom[5][20] = -32'd2683;
    weight_rom[5][21] = -32'd470;
    weight_rom[5][22] = -32'd3556;
    weight_rom[5][23] = 32'd5674;
    weight_rom[5][24] = -32'd5165;
    weight_rom[5][25] = 32'd4429;
    weight_rom[5][26] = -32'd3998;
    weight_rom[5][27] = -32'd4506;
    weight_rom[5][28] = -32'd3979;
    weight_rom[5][29] = -32'd5518;
    weight_rom[5][30] = 32'd2050;
    weight_rom[5][31] = 32'd2745;
    weight_rom[5][32] = -32'd964;
    weight_rom[5][33] = -32'd4064;
    weight_rom[5][34] = 32'd1646;
    weight_rom[5][35] = 32'd3175;
    weight_rom[5][36] = -32'd5124;
    weight_rom[5][37] = -32'd5103;
    weight_rom[5][38] = 32'd4120;
    weight_rom[5][39] = -32'd2256;
    weight_rom[5][40] = 32'd1446;
    weight_rom[5][41] = -32'd5462;
    weight_rom[5][42] = 32'd59;
    weight_rom[5][43] = -32'd472;
    weight_rom[5][44] = 32'd4461;
    weight_rom[5][45] = 32'd3112;
    weight_rom[5][46] = -32'd4032;
    weight_rom[5][47] = 32'd4630;
    weight_rom[5][48] = 32'd5848;
    weight_rom[5][49] = -32'd1775;
    weight_rom[5][50] = 32'd5093;
    weight_rom[5][51] = -32'd6434;
    weight_rom[5][52] = -32'd762;
    weight_rom[5][53] = 32'd662;
    weight_rom[5][54] = 32'd5384;
    weight_rom[5][55] = -32'd1532;
    weight_rom[5][56] = 32'd3273;
    weight_rom[5][57] = -32'd913;
    weight_rom[5][58] = 32'd2172;
    weight_rom[5][59] = 32'd103;
    weight_rom[5][60] = 32'd3513;
    weight_rom[5][61] = -32'd897;
    weight_rom[5][62] = 32'd1848;
    weight_rom[5][63] = 32'd926;
    weight_rom[6][0] = -32'd5792;
    weight_rom[6][1] = 32'd5805;
    weight_rom[6][2] = -32'd4717;
    weight_rom[6][3] = 32'd6429;
    weight_rom[6][4] = 32'd6386;
    weight_rom[6][5] = 32'd1226;
    weight_rom[6][6] = 32'd3896;
    weight_rom[6][7] = -32'd4175;
    weight_rom[6][8] = -32'd6068;
    weight_rom[6][9] = 32'd4873;
    weight_rom[6][10] = -32'd5401;
    weight_rom[6][11] = 32'd408;
    weight_rom[6][12] = 32'd882;
    weight_rom[6][13] = -32'd1564;
    weight_rom[6][14] = -32'd5619;
    weight_rom[6][15] = 32'd1156;
    weight_rom[6][16] = 32'd4587;
    weight_rom[6][17] = -32'd6118;
    weight_rom[6][18] = 32'd97;
    weight_rom[6][19] = 32'd542;
    weight_rom[6][20] = -32'd3507;
    weight_rom[6][21] = 32'd6075;
    weight_rom[6][22] = 32'd1761;
    weight_rom[6][23] = 32'd4292;
    weight_rom[6][24] = -32'd4524;
    weight_rom[6][25] = 32'd4702;
    weight_rom[6][26] = 32'd5117;
    weight_rom[6][27] = 32'd1781;
    weight_rom[6][28] = 32'd5917;
    weight_rom[6][29] = -32'd749;
    weight_rom[6][30] = 32'd6175;
    weight_rom[6][31] = -32'd2995;
    weight_rom[6][32] = 32'd631;
    weight_rom[6][33] = 32'd2644;
    weight_rom[6][34] = 32'd938;
    weight_rom[6][35] = -32'd6223;
    weight_rom[6][36] = -32'd3295;
    weight_rom[6][37] = -32'd6087;
    weight_rom[6][38] = -32'd1545;
    weight_rom[6][39] = 32'd4138;
    weight_rom[6][40] = 32'd608;
    weight_rom[6][41] = 32'd4757;
    weight_rom[6][42] = -32'd3134;
    weight_rom[6][43] = -32'd4806;
    weight_rom[6][44] = -32'd6324;
    weight_rom[6][45] = -32'd3239;
    weight_rom[6][46] = -32'd472;
    weight_rom[6][47] = 32'd4668;
    weight_rom[6][48] = 32'd1045;
    weight_rom[6][49] = 32'd4504;
    weight_rom[6][50] = -32'd2240;
    weight_rom[6][51] = -32'd5565;
    weight_rom[6][52] = -32'd2009;
    weight_rom[6][53] = 32'd4271;
    weight_rom[6][54] = 32'd1511;
    weight_rom[6][55] = 32'd3008;
    weight_rom[6][56] = -32'd5284;
    weight_rom[6][57] = -32'd2952;
    weight_rom[6][58] = -32'd2801;
    weight_rom[6][59] = 32'd374;
    weight_rom[6][60] = 32'd3240;
    weight_rom[6][61] = -32'd3539;
    weight_rom[6][62] = 32'd5259;
    weight_rom[6][63] = -32'd844;
    weight_rom[7][0] = 32'd4799;
    weight_rom[7][1] = -32'd2317;
    weight_rom[7][2] = 32'd240;
    weight_rom[7][3] = -32'd1145;
    weight_rom[7][4] = -32'd4582;
    weight_rom[7][5] = 32'd2347;
    weight_rom[7][6] = -32'd4588;
    weight_rom[7][7] = 32'd1088;
    weight_rom[7][8] = 32'd1261;
    weight_rom[7][9] = -32'd6170;
    weight_rom[7][10] = -32'd1957;
    weight_rom[7][11] = 32'd5722;
    weight_rom[7][12] = -32'd3190;
    weight_rom[7][13] = 32'd4954;
    weight_rom[7][14] = -32'd6394;
    weight_rom[7][15] = -32'd249;
    weight_rom[7][16] = 32'd2215;
    weight_rom[7][17] = -32'd2569;
    weight_rom[7][18] = 32'd4905;
    weight_rom[7][19] = -32'd4533;
    weight_rom[7][20] = -32'd2870;
    weight_rom[7][21] = 32'd249;
    weight_rom[7][22] = -32'd3642;
    weight_rom[7][23] = 32'd2584;
    weight_rom[7][24] = 32'd5829;
    weight_rom[7][25] = 32'd3255;
    weight_rom[7][26] = 32'd3276;
    weight_rom[7][27] = 32'd1301;
    weight_rom[7][28] = -32'd4253;
    weight_rom[7][29] = -32'd3131;
    weight_rom[7][30] = 32'd815;
    weight_rom[7][31] = 32'd5298;
    weight_rom[7][32] = -32'd4264;
    weight_rom[7][33] = 32'd740;
    weight_rom[7][34] = -32'd4130;
    weight_rom[7][35] = -32'd1902;
    weight_rom[7][36] = -32'd2399;
    weight_rom[7][37] = 32'd6479;
    weight_rom[7][38] = -32'd4819;
    weight_rom[7][39] = 32'd1275;
    weight_rom[7][40] = -32'd3280;
    weight_rom[7][41] = -32'd254;
    weight_rom[7][42] = -32'd6434;
    weight_rom[7][43] = 32'd5606;
    weight_rom[7][44] = -32'd5911;
    weight_rom[7][45] = -32'd5671;
    weight_rom[7][46] = -32'd3331;
    weight_rom[7][47] = -32'd5252;
    weight_rom[7][48] = 32'd527;
    weight_rom[7][49] = -32'd3998;
    weight_rom[7][50] = -32'd2430;
    weight_rom[7][51] = -32'd3272;
    weight_rom[7][52] = 32'd3230;
    weight_rom[7][53] = -32'd2575;
    weight_rom[7][54] = -32'd1154;
    weight_rom[7][55] = -32'd6286;
    weight_rom[7][56] = -32'd313;
    weight_rom[7][57] = 32'd5082;
    weight_rom[7][58] = -32'd522;
    weight_rom[7][59] = 32'd4071;
    weight_rom[7][60] = -32'd2468;
    weight_rom[7][61] = 32'd208;
    weight_rom[7][62] = -32'd4405;
    weight_rom[7][63] = -32'd1116;
    weight_rom[8][0] = 32'd1325;
    weight_rom[8][1] = 32'd246;
    weight_rom[8][2] = 32'd4946;
    weight_rom[8][3] = -32'd1677;
    weight_rom[8][4] = 32'd1233;
    weight_rom[8][5] = 32'd3790;
    weight_rom[8][6] = -32'd3548;
    weight_rom[8][7] = -32'd1029;
    weight_rom[8][8] = -32'd3538;
    weight_rom[8][9] = 32'd4270;
    weight_rom[8][10] = -32'd6118;
    weight_rom[8][11] = -32'd6037;
    weight_rom[8][12] = 32'd6067;
    weight_rom[8][13] = 32'd4824;
    weight_rom[8][14] = 32'd5983;
    weight_rom[8][15] = 32'd1865;
    weight_rom[8][16] = -32'd494;
    weight_rom[8][17] = 32'd2007;
    weight_rom[8][18] = -32'd84;
    weight_rom[8][19] = 32'd703;
    weight_rom[8][20] = 32'd3977;
    weight_rom[8][21] = 32'd2327;
    weight_rom[8][22] = -32'd2337;
    weight_rom[8][23] = 32'd2809;
    weight_rom[8][24] = 32'd3100;
    weight_rom[8][25] = -32'd796;
    weight_rom[8][26] = 32'd5350;
    weight_rom[8][27] = -32'd4202;
    weight_rom[8][28] = 32'd887;
    weight_rom[8][29] = -32'd2052;
    weight_rom[8][30] = 32'd2814;
    weight_rom[8][31] = -32'd1642;
    weight_rom[8][32] = -32'd2674;
    weight_rom[8][33] = -32'd1853;
    weight_rom[8][34] = -32'd5772;
    weight_rom[8][35] = 32'd3672;
    weight_rom[8][36] = 32'd4047;
    weight_rom[8][37] = -32'd3503;
    weight_rom[8][38] = -32'd3975;
    weight_rom[8][39] = -32'd1394;
    weight_rom[8][40] = -32'd2054;
    weight_rom[8][41] = -32'd5652;
    weight_rom[8][42] = 32'd1943;
    weight_rom[8][43] = 32'd4819;
    weight_rom[8][44] = 32'd953;
    weight_rom[8][45] = -32'd3040;
    weight_rom[8][46] = 32'd5437;
    weight_rom[8][47] = -32'd5364;
    weight_rom[8][48] = -32'd5893;
    weight_rom[8][49] = 32'd4284;
    weight_rom[8][50] = 32'd158;
    weight_rom[8][51] = 32'd2219;
    weight_rom[8][52] = 32'd5157;
    weight_rom[8][53] = -32'd1330;
    weight_rom[8][54] = 32'd5693;
    weight_rom[8][55] = -32'd3864;
    weight_rom[8][56] = 32'd6444;
    weight_rom[8][57] = -32'd6021;
    weight_rom[8][58] = -32'd4018;
    weight_rom[8][59] = 32'd3087;
    weight_rom[8][60] = -32'd2539;
    weight_rom[8][61] = -32'd3230;
    weight_rom[8][62] = -32'd1554;
    weight_rom[8][63] = 32'd3050;
    weight_rom[9][0] = 32'd2727;
    weight_rom[9][1] = 32'd2661;
    weight_rom[9][2] = 32'd3155;
    weight_rom[9][3] = 32'd3623;
    weight_rom[9][4] = -32'd1561;
    weight_rom[9][5] = -32'd20;
    weight_rom[9][6] = 32'd2913;
    weight_rom[9][7] = 32'd5146;
    weight_rom[9][8] = -32'd4973;
    weight_rom[9][9] = -32'd4864;
    weight_rom[9][10] = -32'd5523;
    weight_rom[9][11] = -32'd4953;
    weight_rom[9][12] = -32'd215;
    weight_rom[9][13] = 32'd4009;
    weight_rom[9][14] = 32'd3113;
    weight_rom[9][15] = -32'd5703;
    weight_rom[9][16] = -32'd1156;
    weight_rom[9][17] = 32'd5744;
    weight_rom[9][18] = 32'd2651;
    weight_rom[9][19] = 32'd546;
    weight_rom[9][20] = 32'd5626;
    weight_rom[9][21] = -32'd2465;
    weight_rom[9][22] = 32'd4561;
    weight_rom[9][23] = -32'd501;
    weight_rom[9][24] = 32'd5019;
    weight_rom[9][25] = 32'd1448;
    weight_rom[9][26] = 32'd3391;
    weight_rom[9][27] = 32'd2688;
    weight_rom[9][28] = 32'd1039;
    weight_rom[9][29] = 32'd4385;
    weight_rom[9][30] = -32'd5656;
    weight_rom[9][31] = 32'd653;
    weight_rom[9][32] = 32'd2147;
    weight_rom[9][33] = 32'd5391;
    weight_rom[9][34] = 32'd1367;
    weight_rom[9][35] = 32'd837;
    weight_rom[9][36] = 32'd4921;
    weight_rom[9][37] = -32'd5848;
    weight_rom[9][38] = -32'd3440;
    weight_rom[9][39] = -32'd348;
    weight_rom[9][40] = 32'd4614;
    weight_rom[9][41] = 32'd651;
    weight_rom[9][42] = 32'd145;
    weight_rom[9][43] = 32'd2721;
    weight_rom[9][44] = 32'd4187;
    weight_rom[9][45] = 32'd5402;
    weight_rom[9][46] = -32'd2157;
    weight_rom[9][47] = -32'd3110;
    weight_rom[9][48] = -32'd5729;
    weight_rom[9][49] = 32'd821;
    weight_rom[9][50] = 32'd5776;
    weight_rom[9][51] = 32'd5089;
    weight_rom[9][52] = 32'd3365;
    weight_rom[9][53] = -32'd2399;
    weight_rom[9][54] = -32'd5918;
    weight_rom[9][55] = -32'd169;
    weight_rom[9][56] = 32'd3544;
    weight_rom[9][57] = 32'd5422;
    weight_rom[9][58] = -32'd3796;
    weight_rom[9][59] = 32'd2146;
    weight_rom[9][60] = 32'd4428;
    weight_rom[9][61] = 32'd5774;
    weight_rom[9][62] = -32'd4707;
    weight_rom[9][63] = 32'd2436;
    weight_rom[10][0] = -32'd6283;
    weight_rom[10][1] = -32'd1787;
    weight_rom[10][2] = 32'd2582;
    weight_rom[10][3] = -32'd2086;
    weight_rom[10][4] = 32'd6159;
    weight_rom[10][5] = -32'd5414;
    weight_rom[10][6] = 32'd2884;
    weight_rom[10][7] = 32'd4160;
    weight_rom[10][8] = -32'd5544;
    weight_rom[10][9] = -32'd2161;
    weight_rom[10][10] = -32'd1351;
    weight_rom[10][11] = -32'd626;
    weight_rom[10][12] = 32'd4010;
    weight_rom[10][13] = 32'd3801;
    weight_rom[10][14] = -32'd1923;
    weight_rom[10][15] = 32'd1048;
    weight_rom[10][16] = 32'd1978;
    weight_rom[10][17] = 32'd4865;
    weight_rom[10][18] = 32'd6459;
    weight_rom[10][19] = 32'd3432;
    weight_rom[10][20] = -32'd1243;
    weight_rom[10][21] = 32'd3591;
    weight_rom[10][22] = 32'd2999;
    weight_rom[10][23] = 32'd5518;
    weight_rom[10][24] = -32'd3897;
    weight_rom[10][25] = -32'd4451;
    weight_rom[10][26] = 32'd1273;
    weight_rom[10][27] = -32'd587;
    weight_rom[10][28] = -32'd135;
    weight_rom[10][29] = 32'd5707;
    weight_rom[10][30] = -32'd1079;
    weight_rom[10][31] = -32'd5890;
    weight_rom[10][32] = 32'd6098;
    weight_rom[10][33] = -32'd6279;
    weight_rom[10][34] = 32'd3456;
    weight_rom[10][35] = -32'd3130;
    weight_rom[10][36] = -32'd2589;
    weight_rom[10][37] = -32'd4064;
    weight_rom[10][38] = -32'd2622;
    weight_rom[10][39] = 32'd4647;
    weight_rom[10][40] = 32'd776;
    weight_rom[10][41] = -32'd1085;
    weight_rom[10][42] = -32'd714;
    weight_rom[10][43] = -32'd5161;
    weight_rom[10][44] = -32'd2270;
    weight_rom[10][45] = 32'd1745;
    weight_rom[10][46] = 32'd5927;
    weight_rom[10][47] = 32'd4912;
    weight_rom[10][48] = -32'd4098;
    weight_rom[10][49] = 32'd3436;
    weight_rom[10][50] = -32'd5927;
    weight_rom[10][51] = -32'd525;
    weight_rom[10][52] = -32'd2202;
    weight_rom[10][53] = -32'd427;
    weight_rom[10][54] = -32'd3797;
    weight_rom[10][55] = 32'd4957;
    weight_rom[10][56] = -32'd3794;
    weight_rom[10][57] = 32'd4364;
    weight_rom[10][58] = -32'd6251;
    weight_rom[10][59] = -32'd5067;
    weight_rom[10][60] = -32'd5605;
    weight_rom[10][61] = 32'd5320;
    weight_rom[10][62] = 32'd1637;
    weight_rom[10][63] = 32'd4368;
    weight_rom[11][0] = 32'd6159;
    weight_rom[11][1] = 32'd6183;
    weight_rom[11][2] = 32'd2654;
    weight_rom[11][3] = 32'd5645;
    weight_rom[11][4] = 32'd4484;
    weight_rom[11][5] = 32'd486;
    weight_rom[11][6] = 32'd1850;
    weight_rom[11][7] = -32'd2073;
    weight_rom[11][8] = 32'd2572;
    weight_rom[11][9] = 32'd3191;
    weight_rom[11][10] = -32'd4814;
    weight_rom[11][11] = 32'd5686;
    weight_rom[11][12] = 32'd658;
    weight_rom[11][13] = -32'd2560;
    weight_rom[11][14] = -32'd2666;
    weight_rom[11][15] = 32'd805;
    weight_rom[11][16] = 32'd595;
    weight_rom[11][17] = 32'd3487;
    weight_rom[11][18] = -32'd4830;
    weight_rom[11][19] = 32'd4373;
    weight_rom[11][20] = 32'd5322;
    weight_rom[11][21] = 32'd3577;
    weight_rom[11][22] = -32'd5303;
    weight_rom[11][23] = 32'd2550;
    weight_rom[11][24] = 32'd1147;
    weight_rom[11][25] = 32'd2275;
    weight_rom[11][26] = 32'd2020;
    weight_rom[11][27] = 32'd2198;
    weight_rom[11][28] = 32'd1897;
    weight_rom[11][29] = -32'd4119;
    weight_rom[11][30] = -32'd5028;
    weight_rom[11][31] = -32'd968;
    weight_rom[11][32] = -32'd5892;
    weight_rom[11][33] = -32'd2414;
    weight_rom[11][34] = 32'd306;
    weight_rom[11][35] = 32'd2555;
    weight_rom[11][36] = 32'd4701;
    weight_rom[11][37] = -32'd6042;
    weight_rom[11][38] = 32'd1871;
    weight_rom[11][39] = -32'd2097;
    weight_rom[11][40] = 32'd193;
    weight_rom[11][41] = 32'd4951;
    weight_rom[11][42] = 32'd6120;
    weight_rom[11][43] = 32'd3615;
    weight_rom[11][44] = -32'd1971;
    weight_rom[11][45] = 32'd2897;
    weight_rom[11][46] = 32'd433;
    weight_rom[11][47] = -32'd4864;
    weight_rom[11][48] = -32'd6128;
    weight_rom[11][49] = 32'd2799;
    weight_rom[11][50] = -32'd1936;
    weight_rom[11][51] = 32'd1402;
    weight_rom[11][52] = 32'd3203;
    weight_rom[11][53] = -32'd2810;
    weight_rom[11][54] = 32'd863;
    weight_rom[11][55] = 32'd357;
    weight_rom[11][56] = 32'd18;
    weight_rom[11][57] = -32'd2653;
    weight_rom[11][58] = 32'd5200;
    weight_rom[11][59] = 32'd2891;
    weight_rom[11][60] = 32'd4995;
    weight_rom[11][61] = 32'd875;
    weight_rom[11][62] = 32'd2999;
    weight_rom[11][63] = -32'd3277;
    weight_rom[12][0] = 32'd4357;
    weight_rom[12][1] = 32'd6061;
    weight_rom[12][2] = -32'd1841;
    weight_rom[12][3] = 32'd4697;
    weight_rom[12][4] = 32'd4434;
    weight_rom[12][5] = 32'd1138;
    weight_rom[12][6] = 32'd2542;
    weight_rom[12][7] = -32'd3153;
    weight_rom[12][8] = -32'd2098;
    weight_rom[12][9] = -32'd4446;
    weight_rom[12][10] = 32'd885;
    weight_rom[12][11] = -32'd2409;
    weight_rom[12][12] = -32'd5984;
    weight_rom[12][13] = -32'd5492;
    weight_rom[12][14] = -32'd1969;
    weight_rom[12][15] = 32'd795;
    weight_rom[12][16] = -32'd5737;
    weight_rom[12][17] = 32'd3780;
    weight_rom[12][18] = -32'd2952;
    weight_rom[12][19] = -32'd780;
    weight_rom[12][20] = -32'd2339;
    weight_rom[12][21] = 32'd279;
    weight_rom[12][22] = -32'd934;
    weight_rom[12][23] = 32'd3001;
    weight_rom[12][24] = 32'd2636;
    weight_rom[12][25] = -32'd4204;
    weight_rom[12][26] = 32'd5100;
    weight_rom[12][27] = 32'd4421;
    weight_rom[12][28] = -32'd3541;
    weight_rom[12][29] = -32'd1671;
    weight_rom[12][30] = 32'd1478;
    weight_rom[12][31] = 32'd4356;
    weight_rom[12][32] = 32'd5116;
    weight_rom[12][33] = -32'd5808;
    weight_rom[12][34] = -32'd3581;
    weight_rom[12][35] = 32'd883;
    weight_rom[12][36] = 32'd4682;
    weight_rom[12][37] = -32'd1418;
    weight_rom[12][38] = 32'd1323;
    weight_rom[12][39] = 32'd4845;
    weight_rom[12][40] = -32'd5248;
    weight_rom[12][41] = -32'd3879;
    weight_rom[12][42] = 32'd933;
    weight_rom[12][43] = 32'd4036;
    weight_rom[12][44] = 32'd1262;
    weight_rom[12][45] = -32'd3183;
    weight_rom[12][46] = 32'd1724;
    weight_rom[12][47] = 32'd2883;
    weight_rom[12][48] = 32'd3189;
    weight_rom[12][49] = -32'd3833;
    weight_rom[12][50] = 32'd4673;
    weight_rom[12][51] = -32'd4082;
    weight_rom[12][52] = -32'd4561;
    weight_rom[12][53] = 32'd6050;
    weight_rom[12][54] = 32'd1514;
    weight_rom[12][55] = 32'd5634;
    weight_rom[12][56] = -32'd3491;
    weight_rom[12][57] = 32'd3791;
    weight_rom[12][58] = -32'd3791;
    weight_rom[12][59] = 32'd3;
    weight_rom[12][60] = -32'd3189;
    weight_rom[12][61] = -32'd1908;
    weight_rom[12][62] = 32'd5661;
    weight_rom[12][63] = 32'd1435;
    weight_rom[13][0] = -32'd3770;
    weight_rom[13][1] = -32'd3253;
    weight_rom[13][2] = -32'd2705;
    weight_rom[13][3] = -32'd930;
    weight_rom[13][4] = -32'd410;
    weight_rom[13][5] = 32'd3217;
    weight_rom[13][6] = 32'd560;
    weight_rom[13][7] = -32'd1576;
    weight_rom[13][8] = 32'd2946;
    weight_rom[13][9] = 32'd4167;
    weight_rom[13][10] = 32'd2483;
    weight_rom[13][11] = 32'd94;
    weight_rom[13][12] = 32'd1745;
    weight_rom[13][13] = -32'd1271;
    weight_rom[13][14] = 32'd3599;
    weight_rom[13][15] = 32'd1356;
    weight_rom[13][16] = 32'd163;
    weight_rom[13][17] = 32'd2162;
    weight_rom[13][18] = -32'd1381;
    weight_rom[13][19] = -32'd2590;
    weight_rom[13][20] = -32'd308;
    weight_rom[13][21] = 32'd6239;
    weight_rom[13][22] = -32'd6171;
    weight_rom[13][23] = 32'd4740;
    weight_rom[13][24] = 32'd2360;
    weight_rom[13][25] = 32'd2542;
    weight_rom[13][26] = 32'd1032;
    weight_rom[13][27] = -32'd4328;
    weight_rom[13][28] = 32'd690;
    weight_rom[13][29] = 32'd5618;
    weight_rom[13][30] = 32'd5747;
    weight_rom[13][31] = 32'd4006;
    weight_rom[13][32] = 32'd1007;
    weight_rom[13][33] = 32'd3493;
    weight_rom[13][34] = 32'd2182;
    weight_rom[13][35] = 32'd3882;
    weight_rom[13][36] = 32'd3468;
    weight_rom[13][37] = 32'd3963;
    weight_rom[13][38] = 32'd2570;
    weight_rom[13][39] = -32'd5398;
    weight_rom[13][40] = -32'd6343;
    weight_rom[13][41] = 32'd4279;
    weight_rom[13][42] = 32'd4763;
    weight_rom[13][43] = 32'd3509;
    weight_rom[13][44] = -32'd2959;
    weight_rom[13][45] = 32'd2875;
    weight_rom[13][46] = 32'd562;
    weight_rom[13][47] = -32'd5227;
    weight_rom[13][48] = 32'd2927;
    weight_rom[13][49] = 32'd901;
    weight_rom[13][50] = -32'd1362;
    weight_rom[13][51] = 32'd3997;
    weight_rom[13][52] = -32'd4845;
    weight_rom[13][53] = -32'd2453;
    weight_rom[13][54] = -32'd6035;
    weight_rom[13][55] = -32'd212;
    weight_rom[13][56] = -32'd1185;
    weight_rom[13][57] = -32'd6144;
    weight_rom[13][58] = -32'd3571;
    weight_rom[13][59] = 32'd5165;
    weight_rom[13][60] = 32'd1218;
    weight_rom[13][61] = -32'd1557;
    weight_rom[13][62] = -32'd2898;
    weight_rom[13][63] = 32'd1116;
    weight_rom[14][0] = -32'd4170;
    weight_rom[14][1] = -32'd36;
    weight_rom[14][2] = 32'd4054;
    weight_rom[14][3] = 32'd3288;
    weight_rom[14][4] = -32'd1116;
    weight_rom[14][5] = -32'd895;
    weight_rom[14][6] = -32'd3253;
    weight_rom[14][7] = 32'd1183;
    weight_rom[14][8] = -32'd5696;
    weight_rom[14][9] = 32'd4353;
    weight_rom[14][10] = 32'd3939;
    weight_rom[14][11] = -32'd6008;
    weight_rom[14][12] = 32'd5916;
    weight_rom[14][13] = -32'd4279;
    weight_rom[14][14] = 32'd2115;
    weight_rom[14][15] = 32'd2313;
    weight_rom[14][16] = 32'd4016;
    weight_rom[14][17] = -32'd3141;
    weight_rom[14][18] = -32'd1024;
    weight_rom[14][19] = -32'd3154;
    weight_rom[14][20] = -32'd3590;
    weight_rom[14][21] = -32'd4907;
    weight_rom[14][22] = -32'd250;
    weight_rom[14][23] = -32'd2961;
    weight_rom[14][24] = -32'd1203;
    weight_rom[14][25] = -32'd3544;
    weight_rom[14][26] = 32'd1735;
    weight_rom[14][27] = -32'd6302;
    weight_rom[14][28] = -32'd1675;
    weight_rom[14][29] = -32'd5743;
    weight_rom[14][30] = 32'd2120;
    weight_rom[14][31] = -32'd3613;
    weight_rom[14][32] = 32'd837;
    weight_rom[14][33] = 32'd2649;
    weight_rom[14][34] = -32'd5503;
    weight_rom[14][35] = 32'd3080;
    weight_rom[14][36] = -32'd4630;
    weight_rom[14][37] = -32'd2080;
    weight_rom[14][38] = -32'd1802;
    weight_rom[14][39] = 32'd3628;
    weight_rom[14][40] = 32'd6077;
    weight_rom[14][41] = 32'd756;
    weight_rom[14][42] = -32'd4725;
    weight_rom[14][43] = -32'd5059;
    weight_rom[14][44] = -32'd6204;
    weight_rom[14][45] = -32'd6185;
    weight_rom[14][46] = -32'd4857;
    weight_rom[14][47] = 32'd1614;
    weight_rom[14][48] = -32'd4770;
    weight_rom[14][49] = 32'd4819;
    weight_rom[14][50] = -32'd3943;
    weight_rom[14][51] = 32'd6125;
    weight_rom[14][52] = -32'd2023;
    weight_rom[14][53] = -32'd5268;
    weight_rom[14][54] = -32'd1270;
    weight_rom[14][55] = -32'd125;
    weight_rom[14][56] = 32'd3671;
    weight_rom[14][57] = 32'd6119;
    weight_rom[14][58] = -32'd2888;
    weight_rom[14][59] = 32'd5503;
    weight_rom[14][60] = 32'd5714;
    weight_rom[14][61] = -32'd1155;
    weight_rom[14][62] = 32'd5900;
    weight_rom[14][63] = -32'd1707;
    weight_rom[15][0] = -32'd4149;
    weight_rom[15][1] = -32'd2609;
    weight_rom[15][2] = 32'd4064;
    weight_rom[15][3] = 32'd3336;
    weight_rom[15][4] = -32'd2970;
    weight_rom[15][5] = -32'd4881;
    weight_rom[15][6] = -32'd2022;
    weight_rom[15][7] = -32'd3040;
    weight_rom[15][8] = -32'd2421;
    weight_rom[15][9] = 32'd97;
    weight_rom[15][10] = -32'd3930;
    weight_rom[15][11] = -32'd4609;
    weight_rom[15][12] = 32'd1331;
    weight_rom[15][13] = 32'd2555;
    weight_rom[15][14] = -32'd4126;
    weight_rom[15][15] = 32'd3997;
    weight_rom[15][16] = -32'd534;
    weight_rom[15][17] = 32'd5337;
    weight_rom[15][18] = -32'd1166;
    weight_rom[15][19] = -32'd4002;
    weight_rom[15][20] = 32'd1841;
    weight_rom[15][21] = -32'd6331;
    weight_rom[15][22] = 32'd2129;
    weight_rom[15][23] = 32'd4024;
    weight_rom[15][24] = -32'd6351;
    weight_rom[15][25] = -32'd5012;
    weight_rom[15][26] = -32'd4502;
    weight_rom[15][27] = 32'd3658;
    weight_rom[15][28] = 32'd2118;
    weight_rom[15][29] = -32'd5343;
    weight_rom[15][30] = -32'd5546;
    weight_rom[15][31] = -32'd3590;
    weight_rom[15][32] = 32'd3;
    weight_rom[15][33] = -32'd2210;
    weight_rom[15][34] = -32'd762;
    weight_rom[15][35] = 32'd1443;
    weight_rom[15][36] = 32'd2494;
    weight_rom[15][37] = -32'd731;
    weight_rom[15][38] = 32'd4246;
    weight_rom[15][39] = 32'd4555;
    weight_rom[15][40] = -32'd1612;
    weight_rom[15][41] = -32'd5837;
    weight_rom[15][42] = 32'd907;
    weight_rom[15][43] = 32'd1886;
    weight_rom[15][44] = 32'd3083;
    weight_rom[15][45] = -32'd1634;
    weight_rom[15][46] = -32'd1627;
    weight_rom[15][47] = -32'd1886;
    weight_rom[15][48] = 32'd4405;
    weight_rom[15][49] = -32'd889;
    weight_rom[15][50] = -32'd985;
    weight_rom[15][51] = -32'd3033;
    weight_rom[15][52] = 32'd4033;
    weight_rom[15][53] = 32'd351;
    weight_rom[15][54] = 32'd1955;
    weight_rom[15][55] = -32'd4984;
    weight_rom[15][56] = 32'd3555;
    weight_rom[15][57] = 32'd348;
    weight_rom[15][58] = -32'd4883;
    weight_rom[15][59] = -32'd5830;
    weight_rom[15][60] = 32'd2334;
    weight_rom[15][61] = 32'd2982;
    weight_rom[15][62] = -32'd5724;
    weight_rom[15][63] = -32'd182;
    weight_rom[16][0] = -32'd2565;
    weight_rom[16][1] = -32'd2820;
    weight_rom[16][2] = 32'd4811;
    weight_rom[16][3] = -32'd5201;
    weight_rom[16][4] = -32'd5814;
    weight_rom[16][5] = -32'd2834;
    weight_rom[16][6] = -32'd4173;
    weight_rom[16][7] = 32'd1627;
    weight_rom[16][8] = 32'd517;
    weight_rom[16][9] = -32'd6469;
    weight_rom[16][10] = -32'd4358;
    weight_rom[16][11] = 32'd6378;
    weight_rom[16][12] = 32'd4183;
    weight_rom[16][13] = -32'd2017;
    weight_rom[16][14] = -32'd4271;
    weight_rom[16][15] = -32'd3017;
    weight_rom[16][16] = -32'd5872;
    weight_rom[16][17] = 32'd2237;
    weight_rom[16][18] = 32'd5342;
    weight_rom[16][19] = -32'd5797;
    weight_rom[16][20] = 32'd6278;
    weight_rom[16][21] = 32'd3541;
    weight_rom[16][22] = -32'd5000;
    weight_rom[16][23] = -32'd3994;
    weight_rom[16][24] = 32'd1086;
    weight_rom[16][25] = -32'd4387;
    weight_rom[16][26] = -32'd341;
    weight_rom[16][27] = 32'd1437;
    weight_rom[16][28] = -32'd4702;
    weight_rom[16][29] = -32'd4419;
    weight_rom[16][30] = -32'd1904;
    weight_rom[16][31] = 32'd4158;
    weight_rom[16][32] = -32'd5644;
    weight_rom[16][33] = 32'd2302;
    weight_rom[16][34] = -32'd4412;
    weight_rom[16][35] = -32'd154;
    weight_rom[16][36] = 32'd5833;
    weight_rom[16][37] = 32'd2301;
    weight_rom[16][38] = -32'd3878;
    weight_rom[16][39] = -32'd4170;
    weight_rom[16][40] = 32'd1352;
    weight_rom[16][41] = 32'd6184;
    weight_rom[16][42] = 32'd4823;
    weight_rom[16][43] = 32'd4382;
    weight_rom[16][44] = 32'd1646;
    weight_rom[16][45] = 32'd1661;
    weight_rom[16][46] = -32'd5254;
    weight_rom[16][47] = 32'd3786;
    weight_rom[16][48] = -32'd4524;
    weight_rom[16][49] = 32'd6115;
    weight_rom[16][50] = -32'd1500;
    weight_rom[16][51] = -32'd67;
    weight_rom[16][52] = -32'd3324;
    weight_rom[16][53] = -32'd5805;
    weight_rom[16][54] = 32'd2596;
    weight_rom[16][55] = 32'd3966;
    weight_rom[16][56] = -32'd3563;
    weight_rom[16][57] = -32'd2578;
    weight_rom[16][58] = 32'd1825;
    weight_rom[16][59] = 32'd4202;
    weight_rom[16][60] = -32'd1121;
    weight_rom[16][61] = -32'd633;
    weight_rom[16][62] = 32'd1350;
    weight_rom[16][63] = -32'd2440;
    weight_rom[17][0] = 32'd324;
    weight_rom[17][1] = -32'd6070;
    weight_rom[17][2] = 32'd5416;
    weight_rom[17][3] = 32'd5276;
    weight_rom[17][4] = 32'd4780;
    weight_rom[17][5] = -32'd1794;
    weight_rom[17][6] = 32'd5353;
    weight_rom[17][7] = -32'd1187;
    weight_rom[17][8] = 32'd3810;
    weight_rom[17][9] = -32'd2791;
    weight_rom[17][10] = -32'd5182;
    weight_rom[17][11] = 32'd6096;
    weight_rom[17][12] = 32'd5035;
    weight_rom[17][13] = 32'd6233;
    weight_rom[17][14] = -32'd5263;
    weight_rom[17][15] = 32'd4260;
    weight_rom[17][16] = 32'd3752;
    weight_rom[17][17] = 32'd792;
    weight_rom[17][18] = 32'd2805;
    weight_rom[17][19] = -32'd2065;
    weight_rom[17][20] = 32'd1356;
    weight_rom[17][21] = 32'd4025;
    weight_rom[17][22] = -32'd2767;
    weight_rom[17][23] = -32'd2027;
    weight_rom[17][24] = -32'd3236;
    weight_rom[17][25] = -32'd6527;
    weight_rom[17][26] = 32'd2836;
    weight_rom[17][27] = 32'd2616;
    weight_rom[17][28] = 32'd928;
    weight_rom[17][29] = 32'd1248;
    weight_rom[17][30] = 32'd664;
    weight_rom[17][31] = 32'd5641;
    weight_rom[17][32] = -32'd5375;
    weight_rom[17][33] = -32'd1364;
    weight_rom[17][34] = -32'd4135;
    weight_rom[17][35] = -32'd4807;
    weight_rom[17][36] = 32'd2392;
    weight_rom[17][37] = 32'd116;
    weight_rom[17][38] = -32'd405;
    weight_rom[17][39] = -32'd912;
    weight_rom[17][40] = -32'd5508;
    weight_rom[17][41] = 32'd165;
    weight_rom[17][42] = 32'd1089;
    weight_rom[17][43] = 32'd1013;
    weight_rom[17][44] = 32'd1058;
    weight_rom[17][45] = -32'd4638;
    weight_rom[17][46] = 32'd1611;
    weight_rom[17][47] = -32'd3490;
    weight_rom[17][48] = -32'd2606;
    weight_rom[17][49] = -32'd626;
    weight_rom[17][50] = 32'd5444;
    weight_rom[17][51] = -32'd5424;
    weight_rom[17][52] = -32'd5724;
    weight_rom[17][53] = -32'd5104;
    weight_rom[17][54] = 32'd1810;
    weight_rom[17][55] = -32'd3316;
    weight_rom[17][56] = 32'd5534;
    weight_rom[17][57] = -32'd1801;
    weight_rom[17][58] = -32'd5568;
    weight_rom[17][59] = -32'd6059;
    weight_rom[17][60] = 32'd2484;
    weight_rom[17][61] = 32'd4675;
    weight_rom[17][62] = -32'd5804;
    weight_rom[17][63] = -32'd4694;
    weight_rom[18][0] = -32'd892;
    weight_rom[18][1] = 32'd1436;
    weight_rom[18][2] = 32'd148;
    weight_rom[18][3] = 32'd68;
    weight_rom[18][4] = 32'd4101;
    weight_rom[18][5] = 32'd1912;
    weight_rom[18][6] = 32'd1093;
    weight_rom[18][7] = 32'd682;
    weight_rom[18][8] = -32'd2375;
    weight_rom[18][9] = 32'd1532;
    weight_rom[18][10] = 32'd1788;
    weight_rom[18][11] = -32'd6488;
    weight_rom[18][12] = -32'd3564;
    weight_rom[18][13] = 32'd1847;
    weight_rom[18][14] = 32'd2101;
    weight_rom[18][15] = -32'd22;
    weight_rom[18][16] = -32'd3914;
    weight_rom[18][17] = -32'd5098;
    weight_rom[18][18] = 32'd1414;
    weight_rom[18][19] = -32'd3011;
    weight_rom[18][20] = -32'd1863;
    weight_rom[18][21] = -32'd4978;
    weight_rom[18][22] = -32'd1339;
    weight_rom[18][23] = -32'd2154;
    weight_rom[18][24] = -32'd652;
    weight_rom[18][25] = 32'd2867;
    weight_rom[18][26] = -32'd3002;
    weight_rom[18][27] = 32'd4432;
    weight_rom[18][28] = -32'd4125;
    weight_rom[18][29] = -32'd4581;
    weight_rom[18][30] = -32'd1268;
    weight_rom[18][31] = -32'd5303;
    weight_rom[18][32] = 32'd1322;
    weight_rom[18][33] = 32'd3358;
    weight_rom[18][34] = -32'd3902;
    weight_rom[18][35] = -32'd3128;
    weight_rom[18][36] = -32'd2207;
    weight_rom[18][37] = 32'd4737;
    weight_rom[18][38] = 32'd3944;
    weight_rom[18][39] = -32'd4384;
    weight_rom[18][40] = 32'd2400;
    weight_rom[18][41] = -32'd2741;
    weight_rom[18][42] = 32'd2857;
    weight_rom[18][43] = 32'd1918;
    weight_rom[18][44] = 32'd3167;
    weight_rom[18][45] = 32'd4233;
    weight_rom[18][46] = -32'd696;
    weight_rom[18][47] = 32'd1824;
    weight_rom[18][48] = -32'd3290;
    weight_rom[18][49] = -32'd4682;
    weight_rom[18][50] = 32'd3433;
    weight_rom[18][51] = 32'd775;
    weight_rom[18][52] = -32'd4827;
    weight_rom[18][53] = -32'd3678;
    weight_rom[18][54] = -32'd2351;
    weight_rom[18][55] = 32'd5237;
    weight_rom[18][56] = 32'd1213;
    weight_rom[18][57] = -32'd5683;
    weight_rom[18][58] = -32'd4794;
    weight_rom[18][59] = -32'd1741;
    weight_rom[18][60] = -32'd2044;
    weight_rom[18][61] = 32'd5820;
    weight_rom[18][62] = 32'd5161;
    weight_rom[18][63] = -32'd3751;
    weight_rom[19][0] = -32'd2736;
    weight_rom[19][1] = 32'd35;
    weight_rom[19][2] = 32'd19;
    weight_rom[19][3] = 32'd4278;
    weight_rom[19][4] = 32'd6549;
    weight_rom[19][5] = 32'd927;
    weight_rom[19][6] = -32'd1299;
    weight_rom[19][7] = -32'd837;
    weight_rom[19][8] = 32'd1650;
    weight_rom[19][9] = 32'd6306;
    weight_rom[19][10] = 32'd2706;
    weight_rom[19][11] = 32'd5921;
    weight_rom[19][12] = -32'd3774;
    weight_rom[19][13] = 32'd4226;
    weight_rom[19][14] = 32'd3465;
    weight_rom[19][15] = -32'd5543;
    weight_rom[19][16] = -32'd3163;
    weight_rom[19][17] = -32'd693;
    weight_rom[19][18] = -32'd2498;
    weight_rom[19][19] = 32'd6113;
    weight_rom[19][20] = 32'd1937;
    weight_rom[19][21] = -32'd3072;
    weight_rom[19][22] = 32'd5498;
    weight_rom[19][23] = 32'd6272;
    weight_rom[19][24] = 32'd5997;
    weight_rom[19][25] = 32'd3046;
    weight_rom[19][26] = -32'd3902;
    weight_rom[19][27] = 32'd3968;
    weight_rom[19][28] = -32'd2901;
    weight_rom[19][29] = 32'd6135;
    weight_rom[19][30] = 32'd4373;
    weight_rom[19][31] = -32'd654;
    weight_rom[19][32] = -32'd2084;
    weight_rom[19][33] = -32'd600;
    weight_rom[19][34] = -32'd1484;
    weight_rom[19][35] = -32'd1060;
    weight_rom[19][36] = 32'd7;
    weight_rom[19][37] = 32'd4797;
    weight_rom[19][38] = -32'd4192;
    weight_rom[19][39] = 32'd2708;
    weight_rom[19][40] = 32'd5669;
    weight_rom[19][41] = -32'd401;
    weight_rom[19][42] = -32'd1677;
    weight_rom[19][43] = -32'd545;
    weight_rom[19][44] = 32'd2296;
    weight_rom[19][45] = -32'd3473;
    weight_rom[19][46] = 32'd3643;
    weight_rom[19][47] = -32'd3464;
    weight_rom[19][48] = -32'd1673;
    weight_rom[19][49] = -32'd1449;
    weight_rom[19][50] = 32'd67;
    weight_rom[19][51] = 32'd36;
    weight_rom[19][52] = 32'd4702;
    weight_rom[19][53] = -32'd467;
    weight_rom[19][54] = -32'd5327;
    weight_rom[19][55] = 32'd5384;
    weight_rom[19][56] = -32'd1573;
    weight_rom[19][57] = 32'd6414;
    weight_rom[19][58] = 32'd1897;
    weight_rom[19][59] = 32'd554;
    weight_rom[19][60] = -32'd2919;
    weight_rom[19][61] = -32'd2150;
    weight_rom[19][62] = 32'd390;
    weight_rom[19][63] = -32'd5170;
    weight_rom[20][0] = 32'd1466;
    weight_rom[20][1] = -32'd5878;
    weight_rom[20][2] = 32'd3909;
    weight_rom[20][3] = -32'd2358;
    weight_rom[20][4] = 32'd6509;
    weight_rom[20][5] = -32'd1886;
    weight_rom[20][6] = -32'd498;
    weight_rom[20][7] = -32'd2693;
    weight_rom[20][8] = 32'd5059;
    weight_rom[20][9] = 32'd1727;
    weight_rom[20][10] = -32'd6139;
    weight_rom[20][11] = 32'd1823;
    weight_rom[20][12] = 32'd1454;
    weight_rom[20][13] = -32'd4816;
    weight_rom[20][14] = -32'd3079;
    weight_rom[20][15] = -32'd5786;
    weight_rom[20][16] = -32'd4394;
    weight_rom[20][17] = -32'd519;
    weight_rom[20][18] = 32'd4243;
    weight_rom[20][19] = 32'd756;
    weight_rom[20][20] = -32'd4942;
    weight_rom[20][21] = -32'd6323;
    weight_rom[20][22] = 32'd6465;
    weight_rom[20][23] = 32'd4673;
    weight_rom[20][24] = -32'd1323;
    weight_rom[20][25] = 32'd195;
    weight_rom[20][26] = -32'd2440;
    weight_rom[20][27] = 32'd6041;
    weight_rom[20][28] = -32'd3686;
    weight_rom[20][29] = -32'd698;
    weight_rom[20][30] = 32'd4124;
    weight_rom[20][31] = -32'd2130;
    weight_rom[20][32] = 32'd5469;
    weight_rom[20][33] = -32'd1149;
    weight_rom[20][34] = -32'd5883;
    weight_rom[20][35] = 32'd1301;
    weight_rom[20][36] = 32'd1910;
    weight_rom[20][37] = -32'd6423;
    weight_rom[20][38] = -32'd5113;
    weight_rom[20][39] = 32'd463;
    weight_rom[20][40] = 32'd991;
    weight_rom[20][41] = 32'd4690;
    weight_rom[20][42] = -32'd5341;
    weight_rom[20][43] = 32'd376;
    weight_rom[20][44] = -32'd3855;
    weight_rom[20][45] = 32'd1995;
    weight_rom[20][46] = -32'd3663;
    weight_rom[20][47] = 32'd2800;
    weight_rom[20][48] = -32'd3215;
    weight_rom[20][49] = 32'd5920;
    weight_rom[20][50] = 32'd6401;
    weight_rom[20][51] = -32'd4660;
    weight_rom[20][52] = 32'd1753;
    weight_rom[20][53] = -32'd874;
    weight_rom[20][54] = -32'd955;
    weight_rom[20][55] = 32'd5810;
    weight_rom[20][56] = 32'd25;
    weight_rom[20][57] = -32'd6038;
    weight_rom[20][58] = -32'd2101;
    weight_rom[20][59] = -32'd4612;
    weight_rom[20][60] = 32'd6510;
    weight_rom[20][61] = 32'd795;
    weight_rom[20][62] = 32'd2219;
    weight_rom[20][63] = 32'd2399;
    weight_rom[21][0] = -32'd4725;
    weight_rom[21][1] = -32'd2901;
    weight_rom[21][2] = 32'd1965;
    weight_rom[21][3] = 32'd5184;
    weight_rom[21][4] = 32'd726;
    weight_rom[21][5] = 32'd6376;
    weight_rom[21][6] = 32'd5862;
    weight_rom[21][7] = 32'd5877;
    weight_rom[21][8] = 32'd1518;
    weight_rom[21][9] = -32'd3148;
    weight_rom[21][10] = 32'd5717;
    weight_rom[21][11] = 32'd4822;
    weight_rom[21][12] = -32'd1166;
    weight_rom[21][13] = 32'd4745;
    weight_rom[21][14] = -32'd6279;
    weight_rom[21][15] = -32'd2172;
    weight_rom[21][16] = -32'd2225;
    weight_rom[21][17] = 32'd4778;
    weight_rom[21][18] = 32'd5964;
    weight_rom[21][19] = -32'd2001;
    weight_rom[21][20] = 32'd5094;
    weight_rom[21][21] = -32'd2709;
    weight_rom[21][22] = -32'd5964;
    weight_rom[21][23] = 32'd2636;
    weight_rom[21][24] = 32'd4453;
    weight_rom[21][25] = -32'd4438;
    weight_rom[21][26] = -32'd3388;
    weight_rom[21][27] = 32'd471;
    weight_rom[21][28] = -32'd4157;
    weight_rom[21][29] = 32'd19;
    weight_rom[21][30] = 32'd1465;
    weight_rom[21][31] = 32'd4858;
    weight_rom[21][32] = -32'd1224;
    weight_rom[21][33] = 32'd5698;
    weight_rom[21][34] = -32'd1339;
    weight_rom[21][35] = 32'd179;
    weight_rom[21][36] = 32'd138;
    weight_rom[21][37] = 32'd3644;
    weight_rom[21][38] = 32'd5029;
    weight_rom[21][39] = 32'd1773;
    weight_rom[21][40] = -32'd4900;
    weight_rom[21][41] = -32'd2557;
    weight_rom[21][42] = -32'd551;
    weight_rom[21][43] = -32'd6103;
    weight_rom[21][44] = -32'd1933;
    weight_rom[21][45] = -32'd1242;
    weight_rom[21][46] = -32'd4396;
    weight_rom[21][47] = 32'd4897;
    weight_rom[21][48] = -32'd144;
    weight_rom[21][49] = -32'd2362;
    weight_rom[21][50] = -32'd455;
    weight_rom[21][51] = -32'd759;
    weight_rom[21][52] = -32'd3234;
    weight_rom[21][53] = 32'd3928;
    weight_rom[21][54] = -32'd4865;
    weight_rom[21][55] = 32'd265;
    weight_rom[21][56] = 32'd1377;
    weight_rom[21][57] = 32'd2030;
    weight_rom[21][58] = 32'd2725;
    weight_rom[21][59] = 32'd3228;
    weight_rom[21][60] = 32'd3287;
    weight_rom[21][61] = -32'd5307;
    weight_rom[21][62] = 32'd4346;
    weight_rom[21][63] = 32'd2106;
    weight_rom[22][0] = -32'd2724;
    weight_rom[22][1] = 32'd5351;
    weight_rom[22][2] = 32'd2647;
    weight_rom[22][3] = -32'd1452;
    weight_rom[22][4] = 32'd3525;
    weight_rom[22][5] = 32'd1386;
    weight_rom[22][6] = -32'd4543;
    weight_rom[22][7] = 32'd3455;
    weight_rom[22][8] = -32'd3500;
    weight_rom[22][9] = 32'd1756;
    weight_rom[22][10] = -32'd5872;
    weight_rom[22][11] = -32'd593;
    weight_rom[22][12] = 32'd4454;
    weight_rom[22][13] = 32'd5541;
    weight_rom[22][14] = -32'd5476;
    weight_rom[22][15] = 32'd3734;
    weight_rom[22][16] = 32'd3365;
    weight_rom[22][17] = 32'd611;
    weight_rom[22][18] = 32'd4210;
    weight_rom[22][19] = 32'd1054;
    weight_rom[22][20] = 32'd40;
    weight_rom[22][21] = 32'd3580;
    weight_rom[22][22] = 32'd3421;
    weight_rom[22][23] = 32'd2976;
    weight_rom[22][24] = -32'd4082;
    weight_rom[22][25] = -32'd5458;
    weight_rom[22][26] = -32'd3736;
    weight_rom[22][27] = -32'd150;
    weight_rom[22][28] = 32'd4269;
    weight_rom[22][29] = -32'd3320;
    weight_rom[22][30] = -32'd1658;
    weight_rom[22][31] = -32'd5458;
    weight_rom[22][32] = -32'd4675;
    weight_rom[22][33] = -32'd3265;
    weight_rom[22][34] = 32'd153;
    weight_rom[22][35] = -32'd2776;
    weight_rom[22][36] = -32'd4981;
    weight_rom[22][37] = -32'd514;
    weight_rom[22][38] = -32'd2058;
    weight_rom[22][39] = -32'd3978;
    weight_rom[22][40] = 32'd1071;
    weight_rom[22][41] = -32'd4028;
    weight_rom[22][42] = -32'd1383;
    weight_rom[22][43] = 32'd1821;
    weight_rom[22][44] = -32'd4900;
    weight_rom[22][45] = 32'd1258;
    weight_rom[22][46] = -32'd1227;
    weight_rom[22][47] = -32'd4891;
    weight_rom[22][48] = -32'd1213;
    weight_rom[22][49] = 32'd4824;
    weight_rom[22][50] = -32'd5790;
    weight_rom[22][51] = -32'd2174;
    weight_rom[22][52] = 32'd724;
    weight_rom[22][53] = 32'd3138;
    weight_rom[22][54] = 32'd5867;
    weight_rom[22][55] = 32'd2321;
    weight_rom[22][56] = 32'd784;
    weight_rom[22][57] = -32'd750;
    weight_rom[22][58] = 32'd752;
    weight_rom[22][59] = -32'd6444;
    weight_rom[22][60] = 32'd1896;
    weight_rom[22][61] = -32'd3925;
    weight_rom[22][62] = -32'd4583;
    weight_rom[22][63] = 32'd5906;
    weight_rom[23][0] = -32'd1751;
    weight_rom[23][1] = -32'd3413;
    weight_rom[23][2] = 32'd3877;
    weight_rom[23][3] = -32'd6411;
    weight_rom[23][4] = 32'd5829;
    weight_rom[23][5] = -32'd3444;
    weight_rom[23][6] = 32'd1130;
    weight_rom[23][7] = -32'd4717;
    weight_rom[23][8] = -32'd6233;
    weight_rom[23][9] = 32'd524;
    weight_rom[23][10] = 32'd541;
    weight_rom[23][11] = 32'd204;
    weight_rom[23][12] = 32'd5243;
    weight_rom[23][13] = -32'd169;
    weight_rom[23][14] = 32'd6132;
    weight_rom[23][15] = 32'd2722;
    weight_rom[23][16] = 32'd254;
    weight_rom[23][17] = -32'd1567;
    weight_rom[23][18] = -32'd6533;
    weight_rom[23][19] = -32'd4729;
    weight_rom[23][20] = -32'd663;
    weight_rom[23][21] = 32'd235;
    weight_rom[23][22] = -32'd1681;
    weight_rom[23][23] = 32'd813;
    weight_rom[23][24] = 32'd2260;
    weight_rom[23][25] = -32'd6302;
    weight_rom[23][26] = -32'd985;
    weight_rom[23][27] = -32'd1286;
    weight_rom[23][28] = -32'd2808;
    weight_rom[23][29] = -32'd380;
    weight_rom[23][30] = -32'd3206;
    weight_rom[23][31] = -32'd3786;
    weight_rom[23][32] = 32'd2814;
    weight_rom[23][33] = -32'd4974;
    weight_rom[23][34] = -32'd218;
    weight_rom[23][35] = -32'd6468;
    weight_rom[23][36] = -32'd2463;
    weight_rom[23][37] = 32'd6407;
    weight_rom[23][38] = 32'd2410;
    weight_rom[23][39] = -32'd3778;
    weight_rom[23][40] = 32'd3491;
    weight_rom[23][41] = -32'd4861;
    weight_rom[23][42] = 32'd4811;
    weight_rom[23][43] = -32'd5486;
    weight_rom[23][44] = -32'd4851;
    weight_rom[23][45] = -32'd5145;
    weight_rom[23][46] = 32'd5591;
    weight_rom[23][47] = 32'd4805;
    weight_rom[23][48] = 32'd6377;
    weight_rom[23][49] = 32'd4997;
    weight_rom[23][50] = -32'd3115;
    weight_rom[23][51] = 32'd286;
    weight_rom[23][52] = 32'd361;
    weight_rom[23][53] = -32'd965;
    weight_rom[23][54] = -32'd325;
    weight_rom[23][55] = 32'd3650;
    weight_rom[23][56] = -32'd178;
    weight_rom[23][57] = 32'd5884;
    weight_rom[23][58] = -32'd3197;
    weight_rom[23][59] = -32'd4343;
    weight_rom[23][60] = -32'd1896;
    weight_rom[23][61] = -32'd1134;
    weight_rom[23][62] = -32'd6047;
    weight_rom[23][63] = 32'd3010;
    weight_rom[24][0] = -32'd575;
    weight_rom[24][1] = -32'd4654;
    weight_rom[24][2] = 32'd5111;
    weight_rom[24][3] = 32'd5313;
    weight_rom[24][4] = 32'd4582;
    weight_rom[24][5] = -32'd5219;
    weight_rom[24][6] = 32'd77;
    weight_rom[24][7] = 32'd4829;
    weight_rom[24][8] = 32'd4850;
    weight_rom[24][9] = 32'd3667;
    weight_rom[24][10] = 32'd2740;
    weight_rom[24][11] = -32'd146;
    weight_rom[24][12] = -32'd1921;
    weight_rom[24][13] = 32'd1392;
    weight_rom[24][14] = -32'd2681;
    weight_rom[24][15] = 32'd3782;
    weight_rom[24][16] = -32'd3868;
    weight_rom[24][17] = 32'd6249;
    weight_rom[24][18] = 32'd1787;
    weight_rom[24][19] = -32'd733;
    weight_rom[24][20] = 32'd1125;
    weight_rom[24][21] = -32'd1991;
    weight_rom[24][22] = -32'd1409;
    weight_rom[24][23] = 32'd5860;
    weight_rom[24][24] = 32'd6252;
    weight_rom[24][25] = -32'd4381;
    weight_rom[24][26] = 32'd5345;
    weight_rom[24][27] = -32'd4539;
    weight_rom[24][28] = 32'd5598;
    weight_rom[24][29] = 32'd2122;
    weight_rom[24][30] = -32'd5165;
    weight_rom[24][31] = 32'd3309;
    weight_rom[24][32] = -32'd2708;
    weight_rom[24][33] = 32'd1108;
    weight_rom[24][34] = -32'd1536;
    weight_rom[24][35] = -32'd49;
    weight_rom[24][36] = 32'd3963;
    weight_rom[24][37] = -32'd219;
    weight_rom[24][38] = -32'd6221;
    weight_rom[24][39] = -32'd6009;
    weight_rom[24][40] = -32'd1226;
    weight_rom[24][41] = -32'd2649;
    weight_rom[24][42] = -32'd3355;
    weight_rom[24][43] = -32'd851;
    weight_rom[24][44] = 32'd2309;
    weight_rom[24][45] = -32'd6331;
    weight_rom[24][46] = 32'd2758;
    weight_rom[24][47] = 32'd1226;
    weight_rom[24][48] = -32'd5820;
    weight_rom[24][49] = -32'd1963;
    weight_rom[24][50] = -32'd837;
    weight_rom[24][51] = 32'd1122;
    weight_rom[24][52] = 32'd2037;
    weight_rom[24][53] = -32'd2179;
    weight_rom[24][54] = -32'd2395;
    weight_rom[24][55] = -32'd4836;
    weight_rom[24][56] = 32'd64;
    weight_rom[24][57] = -32'd3329;
    weight_rom[24][58] = 32'd1976;
    weight_rom[24][59] = 32'd1058;
    weight_rom[24][60] = -32'd5909;
    weight_rom[24][61] = -32'd3850;
    weight_rom[24][62] = 32'd4966;
    weight_rom[24][63] = -32'd5871;
    weight_rom[25][0] = 32'd3737;
    weight_rom[25][1] = -32'd138;
    weight_rom[25][2] = -32'd2123;
    weight_rom[25][3] = -32'd5357;
    weight_rom[25][4] = -32'd3311;
    weight_rom[25][5] = -32'd4550;
    weight_rom[25][6] = 32'd1460;
    weight_rom[25][7] = -32'd164;
    weight_rom[25][8] = -32'd6274;
    weight_rom[25][9] = -32'd5151;
    weight_rom[25][10] = 32'd4862;
    weight_rom[25][11] = 32'd2187;
    weight_rom[25][12] = -32'd3448;
    weight_rom[25][13] = 32'd3470;
    weight_rom[25][14] = 32'd3528;
    weight_rom[25][15] = 32'd226;
    weight_rom[25][16] = 32'd4952;
    weight_rom[25][17] = -32'd5102;
    weight_rom[25][18] = -32'd5883;
    weight_rom[25][19] = 32'd1654;
    weight_rom[25][20] = 32'd1635;
    weight_rom[25][21] = -32'd1681;
    weight_rom[25][22] = 32'd3332;
    weight_rom[25][23] = -32'd49;
    weight_rom[25][24] = -32'd5218;
    weight_rom[25][25] = 32'd5123;
    weight_rom[25][26] = 32'd92;
    weight_rom[25][27] = 32'd951;
    weight_rom[25][28] = 32'd6159;
    weight_rom[25][29] = 32'd3292;
    weight_rom[25][30] = -32'd1901;
    weight_rom[25][31] = -32'd5881;
    weight_rom[25][32] = 32'd333;
    weight_rom[25][33] = 32'd6151;
    weight_rom[25][34] = 32'd4445;
    weight_rom[25][35] = -32'd2809;
    weight_rom[25][36] = 32'd4737;
    weight_rom[25][37] = 32'd6381;
    weight_rom[25][38] = 32'd2490;
    weight_rom[25][39] = -32'd2332;
    weight_rom[25][40] = 32'd4978;
    weight_rom[25][41] = 32'd3670;
    weight_rom[25][42] = 32'd6117;
    weight_rom[25][43] = -32'd2717;
    weight_rom[25][44] = 32'd4700;
    weight_rom[25][45] = 32'd5368;
    weight_rom[25][46] = -32'd1062;
    weight_rom[25][47] = -32'd4887;
    weight_rom[25][48] = -32'd4690;
    weight_rom[25][49] = -32'd5462;
    weight_rom[25][50] = -32'd4497;
    weight_rom[25][51] = -32'd6442;
    weight_rom[25][52] = -32'd3497;
    weight_rom[25][53] = -32'd2405;
    weight_rom[25][54] = 32'd3490;
    weight_rom[25][55] = 32'd1323;
    weight_rom[25][56] = -32'd4241;
    weight_rom[25][57] = 32'd420;
    weight_rom[25][58] = -32'd5029;
    weight_rom[25][59] = 32'd2810;
    weight_rom[25][60] = -32'd6146;
    weight_rom[25][61] = 32'd4935;
    weight_rom[25][62] = -32'd2425;
    weight_rom[25][63] = 32'd5036;
    weight_rom[26][0] = -32'd3936;
    weight_rom[26][1] = 32'd6365;
    weight_rom[26][2] = -32'd1630;
    weight_rom[26][3] = -32'd2368;
    weight_rom[26][4] = -32'd648;
    weight_rom[26][5] = -32'd3329;
    weight_rom[26][6] = -32'd6316;
    weight_rom[26][7] = 32'd5171;
    weight_rom[26][8] = 32'd4911;
    weight_rom[26][9] = 32'd3421;
    weight_rom[26][10] = 32'd2806;
    weight_rom[26][11] = -32'd4723;
    weight_rom[26][12] = 32'd3676;
    weight_rom[26][13] = -32'd4261;
    weight_rom[26][14] = 32'd1634;
    weight_rom[26][15] = -32'd783;
    weight_rom[26][16] = 32'd4975;
    weight_rom[26][17] = -32'd1015;
    weight_rom[26][18] = -32'd3177;
    weight_rom[26][19] = -32'd145;
    weight_rom[26][20] = -32'd5612;
    weight_rom[26][21] = -32'd6535;
    weight_rom[26][22] = 32'd5484;
    weight_rom[26][23] = -32'd1566;
    weight_rom[26][24] = -32'd6444;
    weight_rom[26][25] = -32'd3387;
    weight_rom[26][26] = -32'd4090;
    weight_rom[26][27] = -32'd2922;
    weight_rom[26][28] = 32'd934;
    weight_rom[26][29] = 32'd3327;
    weight_rom[26][30] = -32'd1138;
    weight_rom[26][31] = -32'd97;
    weight_rom[26][32] = 32'd2593;
    weight_rom[26][33] = -32'd1601;
    weight_rom[26][34] = -32'd4648;
    weight_rom[26][35] = 32'd3075;
    weight_rom[26][36] = -32'd4753;
    weight_rom[26][37] = 32'd3336;
    weight_rom[26][38] = -32'd2410;
    weight_rom[26][39] = 32'd783;
    weight_rom[26][40] = 32'd1948;
    weight_rom[26][41] = -32'd371;
    weight_rom[26][42] = 32'd6004;
    weight_rom[26][43] = 32'd595;
    weight_rom[26][44] = 32'd6065;
    weight_rom[26][45] = -32'd3019;
    weight_rom[26][46] = 32'd226;
    weight_rom[26][47] = -32'd949;
    weight_rom[26][48] = -32'd5861;
    weight_rom[26][49] = 32'd2943;
    weight_rom[26][50] = 32'd5866;
    weight_rom[26][51] = 32'd3421;
    weight_rom[26][52] = 32'd4776;
    weight_rom[26][53] = 32'd3591;
    weight_rom[26][54] = -32'd26;
    weight_rom[26][55] = -32'd6104;
    weight_rom[26][56] = 32'd4099;
    weight_rom[26][57] = -32'd231;
    weight_rom[26][58] = 32'd477;
    weight_rom[26][59] = 32'd5461;
    weight_rom[26][60] = 32'd710;
    weight_rom[26][61] = -32'd4478;
    weight_rom[26][62] = -32'd4863;
    weight_rom[26][63] = 32'd4753;
    weight_rom[27][0] = 32'd186;
    weight_rom[27][1] = -32'd3380;
    weight_rom[27][2] = -32'd5321;
    weight_rom[27][3] = 32'd5899;
    weight_rom[27][4] = -32'd4860;
    weight_rom[27][5] = -32'd4447;
    weight_rom[27][6] = 32'd4877;
    weight_rom[27][7] = 32'd3930;
    weight_rom[27][8] = 32'd379;
    weight_rom[27][9] = 32'd540;
    weight_rom[27][10] = 32'd3954;
    weight_rom[27][11] = -32'd6160;
    weight_rom[27][12] = -32'd2951;
    weight_rom[27][13] = 32'd33;
    weight_rom[27][14] = -32'd1547;
    weight_rom[27][15] = -32'd4620;
    weight_rom[27][16] = 32'd4857;
    weight_rom[27][17] = -32'd6002;
    weight_rom[27][18] = -32'd5773;
    weight_rom[27][19] = -32'd1287;
    weight_rom[27][20] = 32'd2393;
    weight_rom[27][21] = -32'd2624;
    weight_rom[27][22] = 32'd5910;
    weight_rom[27][23] = -32'd4416;
    weight_rom[27][24] = -32'd870;
    weight_rom[27][25] = -32'd1910;
    weight_rom[27][26] = -32'd5544;
    weight_rom[27][27] = 32'd5522;
    weight_rom[27][28] = -32'd4679;
    weight_rom[27][29] = 32'd1020;
    weight_rom[27][30] = 32'd2304;
    weight_rom[27][31] = -32'd758;
    weight_rom[27][32] = 32'd5246;
    weight_rom[27][33] = -32'd5740;
    weight_rom[27][34] = 32'd74;
    weight_rom[27][35] = -32'd6239;
    weight_rom[27][36] = 32'd5929;
    weight_rom[27][37] = -32'd3295;
    weight_rom[27][38] = -32'd5823;
    weight_rom[27][39] = 32'd4691;
    weight_rom[27][40] = 32'd5233;
    weight_rom[27][41] = -32'd3571;
    weight_rom[27][42] = -32'd3307;
    weight_rom[27][43] = -32'd4804;
    weight_rom[27][44] = 32'd1682;
    weight_rom[27][45] = 32'd4190;
    weight_rom[27][46] = -32'd5449;
    weight_rom[27][47] = -32'd4445;
    weight_rom[27][48] = 32'd1649;
    weight_rom[27][49] = -32'd2470;
    weight_rom[27][50] = 32'd3497;
    weight_rom[27][51] = 32'd2792;
    weight_rom[27][52] = -32'd2498;
    weight_rom[27][53] = -32'd5871;
    weight_rom[27][54] = -32'd2489;
    weight_rom[27][55] = -32'd31;
    weight_rom[27][56] = 32'd547;
    weight_rom[27][57] = 32'd2658;
    weight_rom[27][58] = -32'd823;
    weight_rom[27][59] = 32'd2693;
    weight_rom[27][60] = 32'd3434;
    weight_rom[27][61] = -32'd581;
    weight_rom[27][62] = -32'd413;
    weight_rom[27][63] = -32'd742;
    weight_rom[28][0] = 32'd1211;
    weight_rom[28][1] = 32'd2256;
    weight_rom[28][2] = 32'd1026;
    weight_rom[28][3] = 32'd5906;
    weight_rom[28][4] = 32'd5951;
    weight_rom[28][5] = -32'd4108;
    weight_rom[28][6] = 32'd5663;
    weight_rom[28][7] = -32'd980;
    weight_rom[28][8] = 32'd5754;
    weight_rom[28][9] = 32'd6068;
    weight_rom[28][10] = -32'd2104;
    weight_rom[28][11] = -32'd2517;
    weight_rom[28][12] = 32'd4228;
    weight_rom[28][13] = -32'd1328;
    weight_rom[28][14] = -32'd3857;
    weight_rom[28][15] = -32'd2251;
    weight_rom[28][16] = -32'd3423;
    weight_rom[28][17] = 32'd3144;
    weight_rom[28][18] = 32'd1360;
    weight_rom[28][19] = 32'd6472;
    weight_rom[28][20] = -32'd3382;
    weight_rom[28][21] = 32'd1919;
    weight_rom[28][22] = 32'd1010;
    weight_rom[28][23] = 32'd3751;
    weight_rom[28][24] = -32'd5339;
    weight_rom[28][25] = -32'd5172;
    weight_rom[28][26] = 32'd2571;
    weight_rom[28][27] = 32'd1090;
    weight_rom[28][28] = -32'd1644;
    weight_rom[28][29] = 32'd5300;
    weight_rom[28][30] = 32'd2073;
    weight_rom[28][31] = -32'd2170;
    weight_rom[28][32] = 32'd3829;
    weight_rom[28][33] = -32'd2106;
    weight_rom[28][34] = -32'd5740;
    weight_rom[28][35] = 32'd1111;
    weight_rom[28][36] = -32'd2243;
    weight_rom[28][37] = 32'd503;
    weight_rom[28][38] = 32'd1439;
    weight_rom[28][39] = 32'd2187;
    weight_rom[28][40] = 32'd1618;
    weight_rom[28][41] = -32'd4375;
    weight_rom[28][42] = -32'd1991;
    weight_rom[28][43] = 32'd2511;
    weight_rom[28][44] = -32'd4140;
    weight_rom[28][45] = 32'd6545;
    weight_rom[28][46] = 32'd6351;
    weight_rom[28][47] = 32'd2626;
    weight_rom[28][48] = -32'd5839;
    weight_rom[28][49] = 32'd3708;
    weight_rom[28][50] = -32'd3037;
    weight_rom[28][51] = -32'd1752;
    weight_rom[28][52] = 32'd2544;
    weight_rom[28][53] = -32'd6385;
    weight_rom[28][54] = 32'd4089;
    weight_rom[28][55] = -32'd4524;
    weight_rom[28][56] = -32'd4835;
    weight_rom[28][57] = -32'd5662;
    weight_rom[28][58] = -32'd3042;
    weight_rom[28][59] = 32'd2251;
    weight_rom[28][60] = 32'd489;
    weight_rom[28][61] = 32'd1385;
    weight_rom[28][62] = 32'd1288;
    weight_rom[28][63] = 32'd1125;
    weight_rom[29][0] = -32'd5944;
    weight_rom[29][1] = 32'd3429;
    weight_rom[29][2] = -32'd6082;
    weight_rom[29][3] = 32'd962;
    weight_rom[29][4] = 32'd1391;
    weight_rom[29][5] = -32'd2816;
    weight_rom[29][6] = 32'd853;
    weight_rom[29][7] = -32'd6259;
    weight_rom[29][8] = 32'd3916;
    weight_rom[29][9] = -32'd2072;
    weight_rom[29][10] = 32'd4126;
    weight_rom[29][11] = 32'd2682;
    weight_rom[29][12] = -32'd999;
    weight_rom[29][13] = -32'd4635;
    weight_rom[29][14] = -32'd4962;
    weight_rom[29][15] = -32'd864;
    weight_rom[29][16] = -32'd639;
    weight_rom[29][17] = 32'd5479;
    weight_rom[29][18] = 32'd2445;
    weight_rom[29][19] = 32'd4984;
    weight_rom[29][20] = 32'd2804;
    weight_rom[29][21] = 32'd6215;
    weight_rom[29][22] = -32'd1872;
    weight_rom[29][23] = 32'd3072;
    weight_rom[29][24] = 32'd3255;
    weight_rom[29][25] = -32'd3639;
    weight_rom[29][26] = -32'd1536;
    weight_rom[29][27] = 32'd1216;
    weight_rom[29][28] = 32'd3902;
    weight_rom[29][29] = 32'd4160;
    weight_rom[29][30] = -32'd5634;
    weight_rom[29][31] = -32'd1381;
    weight_rom[29][32] = 32'd2311;
    weight_rom[29][33] = 32'd77;
    weight_rom[29][34] = -32'd5620;
    weight_rom[29][35] = 32'd5786;
    weight_rom[29][36] = 32'd2127;
    weight_rom[29][37] = 32'd6450;
    weight_rom[29][38] = -32'd3397;
    weight_rom[29][39] = -32'd846;
    weight_rom[29][40] = -32'd4832;
    weight_rom[29][41] = -32'd2192;
    weight_rom[29][42] = 32'd5184;
    weight_rom[29][43] = 32'd3866;
    weight_rom[29][44] = -32'd5168;
    weight_rom[29][45] = -32'd3782;
    weight_rom[29][46] = 32'd2181;
    weight_rom[29][47] = 32'd3393;
    weight_rom[29][48] = 32'd4409;
    weight_rom[29][49] = -32'd751;
    weight_rom[29][50] = 32'd1190;
    weight_rom[29][51] = -32'd5859;
    weight_rom[29][52] = -32'd6342;
    weight_rom[29][53] = 32'd3873;
    weight_rom[29][54] = 32'd4812;
    weight_rom[29][55] = -32'd4155;
    weight_rom[29][56] = 32'd3488;
    weight_rom[29][57] = -32'd4013;
    weight_rom[29][58] = 32'd1363;
    weight_rom[29][59] = -32'd1384;
    weight_rom[29][60] = 32'd4466;
    weight_rom[29][61] = 32'd2514;
    weight_rom[29][62] = -32'd6147;
    weight_rom[29][63] = 32'd6240;
    weight_rom[30][0] = 32'd1409;
    weight_rom[30][1] = -32'd3438;
    weight_rom[30][2] = -32'd450;
    weight_rom[30][3] = 32'd1727;
    weight_rom[30][4] = -32'd3556;
    weight_rom[30][5] = -32'd4281;
    weight_rom[30][6] = 32'd2577;
    weight_rom[30][7] = -32'd3032;
    weight_rom[30][8] = 32'd6526;
    weight_rom[30][9] = 32'd1738;
    weight_rom[30][10] = -32'd5503;
    weight_rom[30][11] = -32'd3907;
    weight_rom[30][12] = 32'd2196;
    weight_rom[30][13] = -32'd1736;
    weight_rom[30][14] = 32'd1507;
    weight_rom[30][15] = -32'd5392;
    weight_rom[30][16] = 32'd6356;
    weight_rom[30][17] = -32'd2883;
    weight_rom[30][18] = -32'd5052;
    weight_rom[30][19] = 32'd1617;
    weight_rom[30][20] = 32'd4227;
    weight_rom[30][21] = 32'd4548;
    weight_rom[30][22] = 32'd3768;
    weight_rom[30][23] = -32'd1515;
    weight_rom[30][24] = 32'd5433;
    weight_rom[30][25] = 32'd251;
    weight_rom[30][26] = 32'd4218;
    weight_rom[30][27] = -32'd1901;
    weight_rom[30][28] = -32'd1738;
    weight_rom[30][29] = 32'd3369;
    weight_rom[30][30] = -32'd1372;
    weight_rom[30][31] = 32'd392;
    weight_rom[30][32] = 32'd2354;
    weight_rom[30][33] = -32'd4431;
    weight_rom[30][34] = 32'd968;
    weight_rom[30][35] = -32'd4267;
    weight_rom[30][36] = 32'd3300;
    weight_rom[30][37] = 32'd4686;
    weight_rom[30][38] = -32'd1483;
    weight_rom[30][39] = 32'd5939;
    weight_rom[30][40] = -32'd2494;
    weight_rom[30][41] = 32'd5766;
    weight_rom[30][42] = 32'd6116;
    weight_rom[30][43] = -32'd4412;
    weight_rom[30][44] = 32'd4100;
    weight_rom[30][45] = -32'd3077;
    weight_rom[30][46] = -32'd2812;
    weight_rom[30][47] = -32'd5166;
    weight_rom[30][48] = 32'd156;
    weight_rom[30][49] = -32'd193;
    weight_rom[30][50] = 32'd2902;
    weight_rom[30][51] = 32'd3341;
    weight_rom[30][52] = -32'd1669;
    weight_rom[30][53] = -32'd299;
    weight_rom[30][54] = 32'd2267;
    weight_rom[30][55] = -32'd1768;
    weight_rom[30][56] = 32'd5668;
    weight_rom[30][57] = -32'd3741;
    weight_rom[30][58] = 32'd4867;
    weight_rom[30][59] = -32'd6536;
    weight_rom[30][60] = -32'd6115;
    weight_rom[30][61] = -32'd1532;
    weight_rom[30][62] = -32'd2950;
    weight_rom[30][63] = 32'd423;
    weight_rom[31][0] = -32'd4318;
    weight_rom[31][1] = 32'd2991;
    weight_rom[31][2] = 32'd558;
    weight_rom[31][3] = -32'd675;
    weight_rom[31][4] = 32'd2250;
    weight_rom[31][5] = 32'd5200;
    weight_rom[31][6] = 32'd5537;
    weight_rom[31][7] = 32'd545;
    weight_rom[31][8] = -32'd1956;
    weight_rom[31][9] = 32'd5662;
    weight_rom[31][10] = 32'd5174;
    weight_rom[31][11] = 32'd2273;
    weight_rom[31][12] = -32'd5301;
    weight_rom[31][13] = -32'd5660;
    weight_rom[31][14] = 32'd3599;
    weight_rom[31][15] = -32'd3662;
    weight_rom[31][16] = 32'd3565;
    weight_rom[31][17] = 32'd4696;
    weight_rom[31][18] = -32'd1522;
    weight_rom[31][19] = 32'd909;
    weight_rom[31][20] = 32'd3984;
    weight_rom[31][21] = -32'd6244;
    weight_rom[31][22] = -32'd3263;
    weight_rom[31][23] = -32'd6223;
    weight_rom[31][24] = -32'd864;
    weight_rom[31][25] = 32'd1412;
    weight_rom[31][26] = 32'd2090;
    weight_rom[31][27] = -32'd5872;
    weight_rom[31][28] = -32'd5413;
    weight_rom[31][29] = -32'd5824;
    weight_rom[31][30] = -32'd4170;
    weight_rom[31][31] = -32'd4438;
    weight_rom[31][32] = 32'd5844;
    weight_rom[31][33] = 32'd2072;
    weight_rom[31][34] = 32'd865;
    weight_rom[31][35] = -32'd371;
    weight_rom[31][36] = 32'd4088;
    weight_rom[31][37] = -32'd5277;
    weight_rom[31][38] = -32'd5497;
    weight_rom[31][39] = 32'd2873;
    weight_rom[31][40] = -32'd3908;
    weight_rom[31][41] = -32'd2057;
    weight_rom[31][42] = -32'd741;
    weight_rom[31][43] = -32'd5186;
    weight_rom[31][44] = 32'd1032;
    weight_rom[31][45] = 32'd2134;
    weight_rom[31][46] = 32'd1124;
    weight_rom[31][47] = 32'd80;
    weight_rom[31][48] = 32'd354;
    weight_rom[31][49] = 32'd3642;
    weight_rom[31][50] = 32'd5783;
    weight_rom[31][51] = 32'd5966;
    weight_rom[31][52] = -32'd1943;
    weight_rom[31][53] = -32'd4838;
    weight_rom[31][54] = -32'd5938;
    weight_rom[31][55] = -32'd885;
    weight_rom[31][56] = 32'd5862;
    weight_rom[31][57] = 32'd3121;
    weight_rom[31][58] = 32'd6539;
    weight_rom[31][59] = -32'd4978;
    weight_rom[31][60] = -32'd1746;
    weight_rom[31][61] = 32'd4837;
    weight_rom[31][62] = -32'd6123;
    weight_rom[31][63] = 32'd5312;
    weight_rom[32][0] = -32'd5700;
    weight_rom[32][1] = -32'd1732;
    weight_rom[32][2] = -32'd2797;
    weight_rom[32][3] = -32'd2710;
    weight_rom[32][4] = 32'd1548;
    weight_rom[32][5] = -32'd5501;
    weight_rom[32][6] = 32'd2716;
    weight_rom[32][7] = 32'd1749;
    weight_rom[32][8] = 32'd3502;
    weight_rom[32][9] = -32'd5209;
    weight_rom[32][10] = 32'd623;
    weight_rom[32][11] = 32'd6159;
    weight_rom[32][12] = 32'd1623;
    weight_rom[32][13] = -32'd6215;
    weight_rom[32][14] = 32'd1886;
    weight_rom[32][15] = 32'd1287;
    weight_rom[32][16] = -32'd6197;
    weight_rom[32][17] = -32'd2723;
    weight_rom[32][18] = -32'd573;
    weight_rom[32][19] = 32'd1581;
    weight_rom[32][20] = 32'd688;
    weight_rom[32][21] = 32'd5224;
    weight_rom[32][22] = 32'd839;
    weight_rom[32][23] = 32'd4443;
    weight_rom[32][24] = -32'd3162;
    weight_rom[32][25] = -32'd3337;
    weight_rom[32][26] = 32'd3882;
    weight_rom[32][27] = -32'd6137;
    weight_rom[32][28] = 32'd744;
    weight_rom[32][29] = -32'd6463;
    weight_rom[32][30] = -32'd4498;
    weight_rom[32][31] = 32'd943;
    weight_rom[32][32] = -32'd2676;
    weight_rom[32][33] = 32'd6524;
    weight_rom[32][34] = 32'd4954;
    weight_rom[32][35] = -32'd5355;
    weight_rom[32][36] = 32'd5842;
    weight_rom[32][37] = 32'd2704;
    weight_rom[32][38] = -32'd4624;
    weight_rom[32][39] = 32'd5638;
    weight_rom[32][40] = 32'd5358;
    weight_rom[32][41] = 32'd6397;
    weight_rom[32][42] = -32'd2346;
    weight_rom[32][43] = -32'd4646;
    weight_rom[32][44] = 32'd1550;
    weight_rom[32][45] = 32'd6100;
    weight_rom[32][46] = -32'd5118;
    weight_rom[32][47] = 32'd4123;
    weight_rom[32][48] = 32'd807;
    weight_rom[32][49] = -32'd1541;
    weight_rom[32][50] = 32'd5002;
    weight_rom[32][51] = -32'd3405;
    weight_rom[32][52] = 32'd569;
    weight_rom[32][53] = -32'd3466;
    weight_rom[32][54] = 32'd869;
    weight_rom[32][55] = 32'd1614;
    weight_rom[32][56] = -32'd1716;
    weight_rom[32][57] = -32'd4074;
    weight_rom[32][58] = 32'd1412;
    weight_rom[32][59] = 32'd452;
    weight_rom[32][60] = -32'd3446;
    weight_rom[32][61] = 32'd895;
    weight_rom[32][62] = -32'd1044;
    weight_rom[32][63] = -32'd5465;
    weight_rom[33][0] = 32'd5883;
    weight_rom[33][1] = 32'd1734;
    weight_rom[33][2] = 32'd1190;
    weight_rom[33][3] = -32'd2245;
    weight_rom[33][4] = -32'd1859;
    weight_rom[33][5] = 32'd321;
    weight_rom[33][6] = -32'd4554;
    weight_rom[33][7] = -32'd3173;
    weight_rom[33][8] = -32'd1285;
    weight_rom[33][9] = 32'd5730;
    weight_rom[33][10] = 32'd4158;
    weight_rom[33][11] = -32'd5322;
    weight_rom[33][12] = -32'd632;
    weight_rom[33][13] = -32'd4781;
    weight_rom[33][14] = 32'd397;
    weight_rom[33][15] = 32'd3088;
    weight_rom[33][16] = -32'd5698;
    weight_rom[33][17] = 32'd5384;
    weight_rom[33][18] = -32'd1716;
    weight_rom[33][19] = -32'd3914;
    weight_rom[33][20] = 32'd264;
    weight_rom[33][21] = 32'd3711;
    weight_rom[33][22] = -32'd1853;
    weight_rom[33][23] = -32'd6403;
    weight_rom[33][24] = -32'd859;
    weight_rom[33][25] = -32'd5796;
    weight_rom[33][26] = -32'd2989;
    weight_rom[33][27] = -32'd1004;
    weight_rom[33][28] = 32'd4523;
    weight_rom[33][29] = -32'd3769;
    weight_rom[33][30] = 32'd4289;
    weight_rom[33][31] = 32'd4003;
    weight_rom[33][32] = -32'd6539;
    weight_rom[33][33] = -32'd632;
    weight_rom[33][34] = 32'd758;
    weight_rom[33][35] = 32'd1647;
    weight_rom[33][36] = -32'd2452;
    weight_rom[33][37] = -32'd2024;
    weight_rom[33][38] = -32'd2647;
    weight_rom[33][39] = 32'd361;
    weight_rom[33][40] = 32'd3413;
    weight_rom[33][41] = -32'd193;
    weight_rom[33][42] = 32'd342;
    weight_rom[33][43] = 32'd4943;
    weight_rom[33][44] = 32'd3689;
    weight_rom[33][45] = 32'd5450;
    weight_rom[33][46] = 32'd6105;
    weight_rom[33][47] = 32'd5716;
    weight_rom[33][48] = -32'd4314;
    weight_rom[33][49] = -32'd745;
    weight_rom[33][50] = 32'd199;
    weight_rom[33][51] = -32'd2313;
    weight_rom[33][52] = -32'd5600;
    weight_rom[33][53] = 32'd5668;
    weight_rom[33][54] = 32'd3451;
    weight_rom[33][55] = -32'd5578;
    weight_rom[33][56] = -32'd4777;
    weight_rom[33][57] = 32'd963;
    weight_rom[33][58] = -32'd1249;
    weight_rom[33][59] = 32'd2295;
    weight_rom[33][60] = -32'd691;
    weight_rom[33][61] = -32'd792;
    weight_rom[33][62] = 32'd5178;
    weight_rom[33][63] = -32'd4049;
    weight_rom[34][0] = 32'd6103;
    weight_rom[34][1] = 32'd1750;
    weight_rom[34][2] = -32'd6153;
    weight_rom[34][3] = 32'd2261;
    weight_rom[34][4] = -32'd5065;
    weight_rom[34][5] = -32'd1174;
    weight_rom[34][6] = 32'd999;
    weight_rom[34][7] = -32'd4727;
    weight_rom[34][8] = -32'd263;
    weight_rom[34][9] = 32'd2462;
    weight_rom[34][10] = -32'd624;
    weight_rom[34][11] = 32'd2262;
    weight_rom[34][12] = 32'd1135;
    weight_rom[34][13] = 32'd6070;
    weight_rom[34][14] = -32'd6003;
    weight_rom[34][15] = 32'd6531;
    weight_rom[34][16] = -32'd472;
    weight_rom[34][17] = 32'd3328;
    weight_rom[34][18] = -32'd4967;
    weight_rom[34][19] = -32'd1374;
    weight_rom[34][20] = -32'd4680;
    weight_rom[34][21] = 32'd3674;
    weight_rom[34][22] = 32'd2052;
    weight_rom[34][23] = 32'd2669;
    weight_rom[34][24] = 32'd2928;
    weight_rom[34][25] = -32'd1428;
    weight_rom[34][26] = 32'd2521;
    weight_rom[34][27] = -32'd5445;
    weight_rom[34][28] = 32'd3878;
    weight_rom[34][29] = 32'd2143;
    weight_rom[34][30] = -32'd6004;
    weight_rom[34][31] = 32'd3409;
    weight_rom[34][32] = -32'd2989;
    weight_rom[34][33] = -32'd1904;
    weight_rom[34][34] = 32'd6026;
    weight_rom[34][35] = 32'd662;
    weight_rom[34][36] = 32'd4698;
    weight_rom[34][37] = -32'd6462;
    weight_rom[34][38] = -32'd5377;
    weight_rom[34][39] = -32'd3160;
    weight_rom[34][40] = 32'd2312;
    weight_rom[34][41] = -32'd4205;
    weight_rom[34][42] = 32'd2461;
    weight_rom[34][43] = 32'd369;
    weight_rom[34][44] = 32'd2664;
    weight_rom[34][45] = 32'd37;
    weight_rom[34][46] = -32'd4262;
    weight_rom[34][47] = 32'd177;
    weight_rom[34][48] = -32'd3962;
    weight_rom[34][49] = -32'd1622;
    weight_rom[34][50] = 32'd3599;
    weight_rom[34][51] = -32'd4144;
    weight_rom[34][52] = 32'd3802;
    weight_rom[34][53] = 32'd4712;
    weight_rom[34][54] = -32'd4764;
    weight_rom[34][55] = 32'd48;
    weight_rom[34][56] = 32'd241;
    weight_rom[34][57] = -32'd3732;
    weight_rom[34][58] = -32'd3601;
    weight_rom[34][59] = -32'd1081;
    weight_rom[34][60] = -32'd5604;
    weight_rom[34][61] = -32'd5672;
    weight_rom[34][62] = 32'd6326;
    weight_rom[34][63] = -32'd776;
    weight_rom[35][0] = 32'd4042;
    weight_rom[35][1] = 32'd468;
    weight_rom[35][2] = -32'd6064;
    weight_rom[35][3] = 32'd3307;
    weight_rom[35][4] = 32'd2248;
    weight_rom[35][5] = 32'd6322;
    weight_rom[35][6] = 32'd1398;
    weight_rom[35][7] = 32'd4389;
    weight_rom[35][8] = 32'd1671;
    weight_rom[35][9] = -32'd5664;
    weight_rom[35][10] = 32'd1881;
    weight_rom[35][11] = -32'd737;
    weight_rom[35][12] = -32'd4351;
    weight_rom[35][13] = 32'd649;
    weight_rom[35][14] = 32'd6140;
    weight_rom[35][15] = 32'd5676;
    weight_rom[35][16] = 32'd5363;
    weight_rom[35][17] = 32'd3996;
    weight_rom[35][18] = -32'd1062;
    weight_rom[35][19] = -32'd6036;
    weight_rom[35][20] = 32'd3609;
    weight_rom[35][21] = -32'd550;
    weight_rom[35][22] = -32'd3402;
    weight_rom[35][23] = 32'd6163;
    weight_rom[35][24] = -32'd6434;
    weight_rom[35][25] = -32'd3483;
    weight_rom[35][26] = -32'd3092;
    weight_rom[35][27] = 32'd1400;
    weight_rom[35][28] = -32'd4258;
    weight_rom[35][29] = -32'd1163;
    weight_rom[35][30] = -32'd1059;
    weight_rom[35][31] = -32'd4536;
    weight_rom[35][32] = -32'd3697;
    weight_rom[35][33] = -32'd1301;
    weight_rom[35][34] = -32'd5915;
    weight_rom[35][35] = -32'd1214;
    weight_rom[35][36] = -32'd4827;
    weight_rom[35][37] = -32'd1265;
    weight_rom[35][38] = 32'd5384;
    weight_rom[35][39] = -32'd5861;
    weight_rom[35][40] = -32'd2608;
    weight_rom[35][41] = 32'd5126;
    weight_rom[35][42] = -32'd2969;
    weight_rom[35][43] = -32'd429;
    weight_rom[35][44] = 32'd4383;
    weight_rom[35][45] = 32'd3868;
    weight_rom[35][46] = 32'd1940;
    weight_rom[35][47] = 32'd5901;
    weight_rom[35][48] = -32'd2374;
    weight_rom[35][49] = -32'd1738;
    weight_rom[35][50] = 32'd814;
    weight_rom[35][51] = 32'd1008;
    weight_rom[35][52] = -32'd3699;
    weight_rom[35][53] = 32'd2749;
    weight_rom[35][54] = -32'd3556;
    weight_rom[35][55] = -32'd4159;
    weight_rom[35][56] = -32'd5077;
    weight_rom[35][57] = 32'd4739;
    weight_rom[35][58] = -32'd3183;
    weight_rom[35][59] = 32'd3023;
    weight_rom[35][60] = 32'd5952;
    weight_rom[35][61] = -32'd462;
    weight_rom[35][62] = 32'd1796;
    weight_rom[35][63] = 32'd1110;
    weight_rom[36][0] = -32'd2560;
    weight_rom[36][1] = -32'd5370;
    weight_rom[36][2] = 32'd4228;
    weight_rom[36][3] = 32'd3821;
    weight_rom[36][4] = 32'd266;
    weight_rom[36][5] = -32'd5085;
    weight_rom[36][6] = -32'd994;
    weight_rom[36][7] = 32'd6349;
    weight_rom[36][8] = 32'd4897;
    weight_rom[36][9] = -32'd2608;
    weight_rom[36][10] = 32'd346;
    weight_rom[36][11] = 32'd4825;
    weight_rom[36][12] = 32'd3104;
    weight_rom[36][13] = 32'd6105;
    weight_rom[36][14] = 32'd3915;
    weight_rom[36][15] = 32'd1868;
    weight_rom[36][16] = 32'd507;
    weight_rom[36][17] = -32'd6317;
    weight_rom[36][18] = 32'd3292;
    weight_rom[36][19] = -32'd320;
    weight_rom[36][20] = -32'd2996;
    weight_rom[36][21] = -32'd1336;
    weight_rom[36][22] = -32'd4042;
    weight_rom[36][23] = -32'd817;
    weight_rom[36][24] = 32'd1172;
    weight_rom[36][25] = -32'd3675;
    weight_rom[36][26] = 32'd5754;
    weight_rom[36][27] = 32'd4993;
    weight_rom[36][28] = 32'd2264;
    weight_rom[36][29] = -32'd1279;
    weight_rom[36][30] = -32'd4348;
    weight_rom[36][31] = -32'd4597;
    weight_rom[36][32] = 32'd2121;
    weight_rom[36][33] = -32'd5044;
    weight_rom[36][34] = -32'd5268;
    weight_rom[36][35] = 32'd280;
    weight_rom[36][36] = 32'd2687;
    weight_rom[36][37] = -32'd3476;
    weight_rom[36][38] = -32'd6474;
    weight_rom[36][39] = 32'd2963;
    weight_rom[36][40] = -32'd4141;
    weight_rom[36][41] = -32'd519;
    weight_rom[36][42] = 32'd3099;
    weight_rom[36][43] = -32'd5154;
    weight_rom[36][44] = -32'd5816;
    weight_rom[36][45] = -32'd4774;
    weight_rom[36][46] = -32'd3336;
    weight_rom[36][47] = 32'd467;
    weight_rom[36][48] = 32'd1225;
    weight_rom[36][49] = 32'd340;
    weight_rom[36][50] = 32'd690;
    weight_rom[36][51] = -32'd4524;
    weight_rom[36][52] = 32'd2320;
    weight_rom[36][53] = -32'd232;
    weight_rom[36][54] = 32'd5013;
    weight_rom[36][55] = 32'd969;
    weight_rom[36][56] = 32'd5688;
    weight_rom[36][57] = 32'd5795;
    weight_rom[36][58] = -32'd269;
    weight_rom[36][59] = 32'd286;
    weight_rom[36][60] = -32'd3627;
    weight_rom[36][61] = 32'd4203;
    weight_rom[36][62] = -32'd4434;
    weight_rom[36][63] = 32'd4144;
    weight_rom[37][0] = -32'd5273;
    weight_rom[37][1] = 32'd4394;
    weight_rom[37][2] = -32'd1832;
    weight_rom[37][3] = 32'd3796;
    weight_rom[37][4] = 32'd3569;
    weight_rom[37][5] = -32'd1338;
    weight_rom[37][6] = 32'd3099;
    weight_rom[37][7] = 32'd336;
    weight_rom[37][8] = 32'd6344;
    weight_rom[37][9] = 32'd2728;
    weight_rom[37][10] = 32'd3035;
    weight_rom[37][11] = -32'd4231;
    weight_rom[37][12] = 32'd4755;
    weight_rom[37][13] = -32'd884;
    weight_rom[37][14] = -32'd2715;
    weight_rom[37][15] = -32'd1032;
    weight_rom[37][16] = -32'd28;
    weight_rom[37][17] = 32'd6066;
    weight_rom[37][18] = -32'd5622;
    weight_rom[37][19] = 32'd563;
    weight_rom[37][20] = -32'd43;
    weight_rom[37][21] = -32'd2583;
    weight_rom[37][22] = 32'd5481;
    weight_rom[37][23] = -32'd3473;
    weight_rom[37][24] = 32'd1484;
    weight_rom[37][25] = 32'd6027;
    weight_rom[37][26] = 32'd1787;
    weight_rom[37][27] = 32'd5018;
    weight_rom[37][28] = -32'd3663;
    weight_rom[37][29] = 32'd5040;
    weight_rom[37][30] = 32'd4971;
    weight_rom[37][31] = -32'd3038;
    weight_rom[37][32] = 32'd1752;
    weight_rom[37][33] = 32'd5023;
    weight_rom[37][34] = -32'd5976;
    weight_rom[37][35] = 32'd5197;
    weight_rom[37][36] = 32'd3171;
    weight_rom[37][37] = 32'd4179;
    weight_rom[37][38] = -32'd211;
    weight_rom[37][39] = -32'd4963;
    weight_rom[37][40] = 32'd3361;
    weight_rom[37][41] = 32'd2748;
    weight_rom[37][42] = -32'd5876;
    weight_rom[37][43] = 32'd1960;
    weight_rom[37][44] = 32'd3244;
    weight_rom[37][45] = 32'd6257;
    weight_rom[37][46] = 32'd2851;
    weight_rom[37][47] = -32'd1386;
    weight_rom[37][48] = -32'd3799;
    weight_rom[37][49] = 32'd4047;
    weight_rom[37][50] = -32'd5049;
    weight_rom[37][51] = -32'd1884;
    weight_rom[37][52] = 32'd3974;
    weight_rom[37][53] = 32'd266;
    weight_rom[37][54] = -32'd6289;
    weight_rom[37][55] = 32'd1800;
    weight_rom[37][56] = -32'd4147;
    weight_rom[37][57] = 32'd242;
    weight_rom[37][58] = -32'd1739;
    weight_rom[37][59] = -32'd5581;
    weight_rom[37][60] = 32'd5535;
    weight_rom[37][61] = 32'd1501;
    weight_rom[37][62] = 32'd5319;
    weight_rom[37][63] = 32'd6399;
    weight_rom[38][0] = 32'd2414;
    weight_rom[38][1] = -32'd2349;
    weight_rom[38][2] = -32'd4888;
    weight_rom[38][3] = -32'd5358;
    weight_rom[38][4] = 32'd264;
    weight_rom[38][5] = 32'd6153;
    weight_rom[38][6] = 32'd5693;
    weight_rom[38][7] = -32'd4303;
    weight_rom[38][8] = 32'd3516;
    weight_rom[38][9] = -32'd5670;
    weight_rom[38][10] = -32'd5483;
    weight_rom[38][11] = 32'd2524;
    weight_rom[38][12] = -32'd3712;
    weight_rom[38][13] = -32'd2466;
    weight_rom[38][14] = 32'd6291;
    weight_rom[38][15] = 32'd1784;
    weight_rom[38][16] = -32'd5171;
    weight_rom[38][17] = 32'd2971;
    weight_rom[38][18] = -32'd5502;
    weight_rom[38][19] = -32'd3568;
    weight_rom[38][20] = -32'd2827;
    weight_rom[38][21] = -32'd5692;
    weight_rom[38][22] = -32'd5219;
    weight_rom[38][23] = 32'd2685;
    weight_rom[38][24] = 32'd1804;
    weight_rom[38][25] = 32'd1524;
    weight_rom[38][26] = -32'd2300;
    weight_rom[38][27] = 32'd2084;
    weight_rom[38][28] = -32'd3693;
    weight_rom[38][29] = 32'd5184;
    weight_rom[38][30] = 32'd747;
    weight_rom[38][31] = -32'd1820;
    weight_rom[38][32] = 32'd1224;
    weight_rom[38][33] = -32'd1116;
    weight_rom[38][34] = -32'd4125;
    weight_rom[38][35] = -32'd3980;
    weight_rom[38][36] = 32'd2329;
    weight_rom[38][37] = -32'd2132;
    weight_rom[38][38] = -32'd4938;
    weight_rom[38][39] = -32'd2585;
    weight_rom[38][40] = -32'd338;
    weight_rom[38][41] = 32'd6340;
    weight_rom[38][42] = -32'd5907;
    weight_rom[38][43] = 32'd4823;
    weight_rom[38][44] = 32'd4598;
    weight_rom[38][45] = 32'd6086;
    weight_rom[38][46] = 32'd3628;
    weight_rom[38][47] = 32'd4563;
    weight_rom[38][48] = -32'd5028;
    weight_rom[38][49] = -32'd1811;
    weight_rom[38][50] = -32'd4900;
    weight_rom[38][51] = 32'd2582;
    weight_rom[38][52] = 32'd811;
    weight_rom[38][53] = 32'd6229;
    weight_rom[38][54] = 32'd3312;
    weight_rom[38][55] = 32'd743;
    weight_rom[38][56] = -32'd3240;
    weight_rom[38][57] = -32'd1935;
    weight_rom[38][58] = 32'd5423;
    weight_rom[38][59] = -32'd4036;
    weight_rom[38][60] = -32'd971;
    weight_rom[38][61] = 32'd4353;
    weight_rom[38][62] = 32'd212;
    weight_rom[38][63] = -32'd1456;
    weight_rom[39][0] = -32'd784;
    weight_rom[39][1] = -32'd4108;
    weight_rom[39][2] = 32'd291;
    weight_rom[39][3] = -32'd73;
    weight_rom[39][4] = 32'd4616;
    weight_rom[39][5] = 32'd4790;
    weight_rom[39][6] = 32'd5578;
    weight_rom[39][7] = -32'd2984;
    weight_rom[39][8] = -32'd1077;
    weight_rom[39][9] = 32'd1077;
    weight_rom[39][10] = -32'd5762;
    weight_rom[39][11] = 32'd4431;
    weight_rom[39][12] = -32'd5299;
    weight_rom[39][13] = 32'd80;
    weight_rom[39][14] = 32'd1335;
    weight_rom[39][15] = 32'd3744;
    weight_rom[39][16] = 32'd2054;
    weight_rom[39][17] = -32'd2559;
    weight_rom[39][18] = -32'd1903;
    weight_rom[39][19] = 32'd6082;
    weight_rom[39][20] = -32'd4799;
    weight_rom[39][21] = -32'd3562;
    weight_rom[39][22] = 32'd78;
    weight_rom[39][23] = 32'd4156;
    weight_rom[39][24] = -32'd3381;
    weight_rom[39][25] = 32'd745;
    weight_rom[39][26] = -32'd3021;
    weight_rom[39][27] = -32'd3784;
    weight_rom[39][28] = 32'd4903;
    weight_rom[39][29] = 32'd5363;
    weight_rom[39][30] = -32'd3520;
    weight_rom[39][31] = -32'd1199;
    weight_rom[39][32] = -32'd6340;
    weight_rom[39][33] = -32'd1477;
    weight_rom[39][34] = 32'd540;
    weight_rom[39][35] = -32'd6257;
    weight_rom[39][36] = -32'd3246;
    weight_rom[39][37] = 32'd4292;
    weight_rom[39][38] = -32'd2520;
    weight_rom[39][39] = 32'd425;
    weight_rom[39][40] = -32'd3594;
    weight_rom[39][41] = -32'd5895;
    weight_rom[39][42] = -32'd1490;
    weight_rom[39][43] = 32'd4301;
    weight_rom[39][44] = -32'd2803;
    weight_rom[39][45] = -32'd4407;
    weight_rom[39][46] = 32'd2273;
    weight_rom[39][47] = -32'd91;
    weight_rom[39][48] = 32'd6161;
    weight_rom[39][49] = 32'd317;
    weight_rom[39][50] = 32'd387;
    weight_rom[39][51] = 32'd787;
    weight_rom[39][52] = 32'd3157;
    weight_rom[39][53] = 32'd6104;
    weight_rom[39][54] = -32'd343;
    weight_rom[39][55] = 32'd3123;
    weight_rom[39][56] = -32'd1223;
    weight_rom[39][57] = -32'd3485;
    weight_rom[39][58] = -32'd1726;
    weight_rom[39][59] = 32'd4456;
    weight_rom[39][60] = 32'd6363;
    weight_rom[39][61] = -32'd78;
    weight_rom[39][62] = -32'd4538;
    weight_rom[39][63] = -32'd5932;
    weight_rom[40][0] = -32'd4953;
    weight_rom[40][1] = -32'd6019;
    weight_rom[40][2] = 32'd3538;
    weight_rom[40][3] = -32'd5799;
    weight_rom[40][4] = 32'd680;
    weight_rom[40][5] = 32'd4155;
    weight_rom[40][6] = -32'd644;
    weight_rom[40][7] = -32'd6312;
    weight_rom[40][8] = -32'd1030;
    weight_rom[40][9] = -32'd2020;
    weight_rom[40][10] = -32'd3314;
    weight_rom[40][11] = 32'd5827;
    weight_rom[40][12] = -32'd6243;
    weight_rom[40][13] = -32'd792;
    weight_rom[40][14] = 32'd1080;
    weight_rom[40][15] = -32'd5002;
    weight_rom[40][16] = 32'd4221;
    weight_rom[40][17] = 32'd4317;
    weight_rom[40][18] = 32'd5789;
    weight_rom[40][19] = 32'd5366;
    weight_rom[40][20] = 32'd1698;
    weight_rom[40][21] = -32'd3321;
    weight_rom[40][22] = -32'd3658;
    weight_rom[40][23] = 32'd608;
    weight_rom[40][24] = 32'd2805;
    weight_rom[40][25] = -32'd1103;
    weight_rom[40][26] = -32'd4051;
    weight_rom[40][27] = 32'd4757;
    weight_rom[40][28] = -32'd3281;
    weight_rom[40][29] = -32'd2439;
    weight_rom[40][30] = 32'd31;
    weight_rom[40][31] = 32'd2355;
    weight_rom[40][32] = 32'd2998;
    weight_rom[40][33] = 32'd2093;
    weight_rom[40][34] = 32'd1908;
    weight_rom[40][35] = 32'd4740;
    weight_rom[40][36] = 32'd4889;
    weight_rom[40][37] = -32'd6545;
    weight_rom[40][38] = 32'd5584;
    weight_rom[40][39] = 32'd844;
    weight_rom[40][40] = 32'd1528;
    weight_rom[40][41] = -32'd5286;
    weight_rom[40][42] = -32'd1920;
    weight_rom[40][43] = 32'd1652;
    weight_rom[40][44] = 32'd1840;
    weight_rom[40][45] = -32'd2628;
    weight_rom[40][46] = 32'd1500;
    weight_rom[40][47] = -32'd368;
    weight_rom[40][48] = -32'd6265;
    weight_rom[40][49] = 32'd2237;
    weight_rom[40][50] = -32'd3029;
    weight_rom[40][51] = -32'd1488;
    weight_rom[40][52] = 32'd2121;
    weight_rom[40][53] = -32'd3732;
    weight_rom[40][54] = -32'd697;
    weight_rom[40][55] = -32'd2154;
    weight_rom[40][56] = -32'd1531;
    weight_rom[40][57] = -32'd5901;
    weight_rom[40][58] = -32'd1658;
    weight_rom[40][59] = 32'd2948;
    weight_rom[40][60] = 32'd708;
    weight_rom[40][61] = -32'd5000;
    weight_rom[40][62] = 32'd5527;
    weight_rom[40][63] = 32'd3947;
    weight_rom[41][0] = -32'd63;
    weight_rom[41][1] = 32'd1191;
    weight_rom[41][2] = -32'd3724;
    weight_rom[41][3] = 32'd649;
    weight_rom[41][4] = 32'd798;
    weight_rom[41][5] = -32'd3173;
    weight_rom[41][6] = -32'd5069;
    weight_rom[41][7] = 32'd5430;
    weight_rom[41][8] = 32'd3114;
    weight_rom[41][9] = 32'd1584;
    weight_rom[41][10] = -32'd4462;
    weight_rom[41][11] = 32'd2401;
    weight_rom[41][12] = 32'd1860;
    weight_rom[41][13] = -32'd5168;
    weight_rom[41][14] = 32'd3251;
    weight_rom[41][15] = -32'd1180;
    weight_rom[41][16] = -32'd1567;
    weight_rom[41][17] = -32'd2863;
    weight_rom[41][18] = 32'd2209;
    weight_rom[41][19] = 32'd2911;
    weight_rom[41][20] = -32'd5841;
    weight_rom[41][21] = -32'd208;
    weight_rom[41][22] = -32'd6043;
    weight_rom[41][23] = 32'd6121;
    weight_rom[41][24] = -32'd5355;
    weight_rom[41][25] = -32'd931;
    weight_rom[41][26] = 32'd2551;
    weight_rom[41][27] = 32'd5060;
    weight_rom[41][28] = -32'd3103;
    weight_rom[41][29] = 32'd2504;
    weight_rom[41][30] = 32'd3034;
    weight_rom[41][31] = -32'd5810;
    weight_rom[41][32] = -32'd2313;
    weight_rom[41][33] = -32'd759;
    weight_rom[41][34] = -32'd5956;
    weight_rom[41][35] = 32'd1010;
    weight_rom[41][36] = -32'd4340;
    weight_rom[41][37] = -32'd2518;
    weight_rom[41][38] = -32'd4434;
    weight_rom[41][39] = 32'd1318;
    weight_rom[41][40] = -32'd6024;
    weight_rom[41][41] = 32'd2889;
    weight_rom[41][42] = -32'd2416;
    weight_rom[41][43] = -32'd5566;
    weight_rom[41][44] = -32'd2435;
    weight_rom[41][45] = -32'd5240;
    weight_rom[41][46] = 32'd5144;
    weight_rom[41][47] = -32'd127;
    weight_rom[41][48] = 32'd3967;
    weight_rom[41][49] = -32'd3021;
    weight_rom[41][50] = -32'd6277;
    weight_rom[41][51] = -32'd1045;
    weight_rom[41][52] = -32'd1893;
    weight_rom[41][53] = 32'd4077;
    weight_rom[41][54] = -32'd6460;
    weight_rom[41][55] = 32'd3474;
    weight_rom[41][56] = 32'd3862;
    weight_rom[41][57] = -32'd3034;
    weight_rom[41][58] = -32'd1526;
    weight_rom[41][59] = 32'd5174;
    weight_rom[41][60] = 32'd5647;
    weight_rom[41][61] = -32'd6374;
    weight_rom[41][62] = 32'd3374;
    weight_rom[41][63] = 32'd1368;
    weight_rom[42][0] = -32'd6102;
    weight_rom[42][1] = 32'd2327;
    weight_rom[42][2] = 32'd1610;
    weight_rom[42][3] = -32'd766;
    weight_rom[42][4] = 32'd4936;
    weight_rom[42][5] = -32'd4313;
    weight_rom[42][6] = 32'd6354;
    weight_rom[42][7] = -32'd5010;
    weight_rom[42][8] = -32'd3423;
    weight_rom[42][9] = -32'd5954;
    weight_rom[42][10] = 32'd4873;
    weight_rom[42][11] = -32'd37;
    weight_rom[42][12] = 32'd1403;
    weight_rom[42][13] = 32'd1845;
    weight_rom[42][14] = 32'd4086;
    weight_rom[42][15] = 32'd4453;
    weight_rom[42][16] = 32'd3612;
    weight_rom[42][17] = 32'd4885;
    weight_rom[42][18] = 32'd2341;
    weight_rom[42][19] = 32'd437;
    weight_rom[42][20] = 32'd3259;
    weight_rom[42][21] = 32'd3243;
    weight_rom[42][22] = -32'd6081;
    weight_rom[42][23] = -32'd5876;
    weight_rom[42][24] = -32'd3941;
    weight_rom[42][25] = 32'd536;
    weight_rom[42][26] = -32'd3686;
    weight_rom[42][27] = -32'd3976;
    weight_rom[42][28] = -32'd6545;
    weight_rom[42][29] = -32'd2993;
    weight_rom[42][30] = 32'd6004;
    weight_rom[42][31] = -32'd6099;
    weight_rom[42][32] = 32'd2163;
    weight_rom[42][33] = 32'd1942;
    weight_rom[42][34] = 32'd5845;
    weight_rom[42][35] = 32'd5120;
    weight_rom[42][36] = -32'd5850;
    weight_rom[42][37] = -32'd3392;
    weight_rom[42][38] = 32'd6105;
    weight_rom[42][39] = -32'd4374;
    weight_rom[42][40] = -32'd2278;
    weight_rom[42][41] = -32'd2859;
    weight_rom[42][42] = -32'd117;
    weight_rom[42][43] = -32'd5080;
    weight_rom[42][44] = 32'd6002;
    weight_rom[42][45] = -32'd2992;
    weight_rom[42][46] = -32'd5523;
    weight_rom[42][47] = 32'd4545;
    weight_rom[42][48] = 32'd3775;
    weight_rom[42][49] = -32'd2916;
    weight_rom[42][50] = 32'd2920;
    weight_rom[42][51] = 32'd814;
    weight_rom[42][52] = 32'd4048;
    weight_rom[42][53] = -32'd3968;
    weight_rom[42][54] = 32'd4186;
    weight_rom[42][55] = -32'd881;
    weight_rom[42][56] = -32'd572;
    weight_rom[42][57] = 32'd2021;
    weight_rom[42][58] = 32'd4412;
    weight_rom[42][59] = -32'd5012;
    weight_rom[42][60] = -32'd6483;
    weight_rom[42][61] = -32'd2579;
    weight_rom[42][62] = 32'd3037;
    weight_rom[42][63] = -32'd3951;
    weight_rom[43][0] = 32'd5365;
    weight_rom[43][1] = -32'd6336;
    weight_rom[43][2] = -32'd5434;
    weight_rom[43][3] = 32'd5081;
    weight_rom[43][4] = -32'd1265;
    weight_rom[43][5] = 32'd2210;
    weight_rom[43][6] = 32'd4442;
    weight_rom[43][7] = 32'd1002;
    weight_rom[43][8] = -32'd5105;
    weight_rom[43][9] = 32'd4869;
    weight_rom[43][10] = -32'd3680;
    weight_rom[43][11] = 32'd1544;
    weight_rom[43][12] = 32'd612;
    weight_rom[43][13] = -32'd3721;
    weight_rom[43][14] = 32'd2051;
    weight_rom[43][15] = -32'd1522;
    weight_rom[43][16] = 32'd6087;
    weight_rom[43][17] = -32'd5077;
    weight_rom[43][18] = -32'd1809;
    weight_rom[43][19] = 32'd4849;
    weight_rom[43][20] = -32'd2390;
    weight_rom[43][21] = -32'd343;
    weight_rom[43][22] = -32'd4256;
    weight_rom[43][23] = 32'd62;
    weight_rom[43][24] = 32'd4947;
    weight_rom[43][25] = 32'd2574;
    weight_rom[43][26] = 32'd1249;
    weight_rom[43][27] = 32'd3111;
    weight_rom[43][28] = 32'd4858;
    weight_rom[43][29] = -32'd4055;
    weight_rom[43][30] = -32'd3664;
    weight_rom[43][31] = -32'd1416;
    weight_rom[43][32] = 32'd741;
    weight_rom[43][33] = -32'd5748;
    weight_rom[43][34] = 32'd4484;
    weight_rom[43][35] = 32'd1270;
    weight_rom[43][36] = 32'd2850;
    weight_rom[43][37] = -32'd3492;
    weight_rom[43][38] = -32'd3856;
    weight_rom[43][39] = -32'd1576;
    weight_rom[43][40] = -32'd412;
    weight_rom[43][41] = -32'd4137;
    weight_rom[43][42] = -32'd2349;
    weight_rom[43][43] = -32'd5907;
    weight_rom[43][44] = -32'd6115;
    weight_rom[43][45] = 32'd4141;
    weight_rom[43][46] = -32'd2216;
    weight_rom[43][47] = 32'd4350;
    weight_rom[43][48] = -32'd2657;
    weight_rom[43][49] = 32'd5680;
    weight_rom[43][50] = -32'd6127;
    weight_rom[43][51] = -32'd6476;
    weight_rom[43][52] = -32'd2690;
    weight_rom[43][53] = -32'd3754;
    weight_rom[43][54] = -32'd1837;
    weight_rom[43][55] = -32'd207;
    weight_rom[43][56] = -32'd4315;
    weight_rom[43][57] = 32'd440;
    weight_rom[43][58] = 32'd1976;
    weight_rom[43][59] = 32'd6425;
    weight_rom[43][60] = 32'd3253;
    weight_rom[43][61] = 32'd2595;
    weight_rom[43][62] = 32'd2741;
    weight_rom[43][63] = -32'd67;
    weight_rom[44][0] = -32'd3161;
    weight_rom[44][1] = 32'd158;
    weight_rom[44][2] = -32'd5876;
    weight_rom[44][3] = -32'd1954;
    weight_rom[44][4] = -32'd4797;
    weight_rom[44][5] = 32'd5627;
    weight_rom[44][6] = -32'd4919;
    weight_rom[44][7] = -32'd2961;
    weight_rom[44][8] = -32'd1905;
    weight_rom[44][9] = 32'd6206;
    weight_rom[44][10] = 32'd6237;
    weight_rom[44][11] = 32'd4835;
    weight_rom[44][12] = -32'd3513;
    weight_rom[44][13] = 32'd1567;
    weight_rom[44][14] = -32'd4874;
    weight_rom[44][15] = 32'd942;
    weight_rom[44][16] = -32'd3882;
    weight_rom[44][17] = 32'd2669;
    weight_rom[44][18] = 32'd1227;
    weight_rom[44][19] = -32'd4841;
    weight_rom[44][20] = -32'd6551;
    weight_rom[44][21] = -32'd5795;
    weight_rom[44][22] = 32'd4807;
    weight_rom[44][23] = 32'd2863;
    weight_rom[44][24] = 32'd3129;
    weight_rom[44][25] = 32'd2649;
    weight_rom[44][26] = -32'd3084;
    weight_rom[44][27] = -32'd2798;
    weight_rom[44][28] = 32'd3835;
    weight_rom[44][29] = -32'd4133;
    weight_rom[44][30] = 32'd5061;
    weight_rom[44][31] = 32'd2584;
    weight_rom[44][32] = -32'd2061;
    weight_rom[44][33] = 32'd4112;
    weight_rom[44][34] = -32'd2665;
    weight_rom[44][35] = 32'd4065;
    weight_rom[44][36] = -32'd321;
    weight_rom[44][37] = -32'd5659;
    weight_rom[44][38] = 32'd3166;
    weight_rom[44][39] = 32'd1536;
    weight_rom[44][40] = -32'd4614;
    weight_rom[44][41] = -32'd6037;
    weight_rom[44][42] = -32'd4033;
    weight_rom[44][43] = -32'd3178;
    weight_rom[44][44] = 32'd1045;
    weight_rom[44][45] = -32'd1594;
    weight_rom[44][46] = -32'd3299;
    weight_rom[44][47] = -32'd1264;
    weight_rom[44][48] = -32'd4775;
    weight_rom[44][49] = 32'd2929;
    weight_rom[44][50] = 32'd1248;
    weight_rom[44][51] = -32'd5524;
    weight_rom[44][52] = 32'd933;
    weight_rom[44][53] = 32'd2308;
    weight_rom[44][54] = 32'd534;
    weight_rom[44][55] = 32'd1941;
    weight_rom[44][56] = -32'd3051;
    weight_rom[44][57] = 32'd5820;
    weight_rom[44][58] = 32'd1496;
    weight_rom[44][59] = -32'd3808;
    weight_rom[44][60] = 32'd5282;
    weight_rom[44][61] = 32'd3804;
    weight_rom[44][62] = -32'd3927;
    weight_rom[44][63] = 32'd3176;
    weight_rom[45][0] = 32'd2130;
    weight_rom[45][1] = -32'd3584;
    weight_rom[45][2] = 32'd410;
    weight_rom[45][3] = -32'd5019;
    weight_rom[45][4] = -32'd6176;
    weight_rom[45][5] = 32'd744;
    weight_rom[45][6] = 32'd5516;
    weight_rom[45][7] = 32'd710;
    weight_rom[45][8] = -32'd2788;
    weight_rom[45][9] = 32'd6145;
    weight_rom[45][10] = -32'd2137;
    weight_rom[45][11] = 32'd925;
    weight_rom[45][12] = -32'd1429;
    weight_rom[45][13] = 32'd1968;
    weight_rom[45][14] = -32'd2119;
    weight_rom[45][15] = 32'd1150;
    weight_rom[45][16] = 32'd305;
    weight_rom[45][17] = 32'd533;
    weight_rom[45][18] = -32'd6420;
    weight_rom[45][19] = 32'd3807;
    weight_rom[45][20] = 32'd145;
    weight_rom[45][21] = 32'd6000;
    weight_rom[45][22] = -32'd2851;
    weight_rom[45][23] = 32'd4753;
    weight_rom[45][24] = -32'd6373;
    weight_rom[45][25] = -32'd4303;
    weight_rom[45][26] = 32'd2122;
    weight_rom[45][27] = 32'd3966;
    weight_rom[45][28] = 32'd1668;
    weight_rom[45][29] = -32'd2069;
    weight_rom[45][30] = 32'd5692;
    weight_rom[45][31] = -32'd4018;
    weight_rom[45][32] = -32'd4789;
    weight_rom[45][33] = 32'd5773;
    weight_rom[45][34] = -32'd5541;
    weight_rom[45][35] = -32'd921;
    weight_rom[45][36] = 32'd4575;
    weight_rom[45][37] = -32'd4100;
    weight_rom[45][38] = 32'd611;
    weight_rom[45][39] = 32'd6158;
    weight_rom[45][40] = 32'd6352;
    weight_rom[45][41] = -32'd6267;
    weight_rom[45][42] = -32'd2497;
    weight_rom[45][43] = -32'd4775;
    weight_rom[45][44] = -32'd4371;
    weight_rom[45][45] = -32'd5394;
    weight_rom[45][46] = 32'd6396;
    weight_rom[45][47] = -32'd2184;
    weight_rom[45][48] = -32'd4644;
    weight_rom[45][49] = 32'd1011;
    weight_rom[45][50] = 32'd513;
    weight_rom[45][51] = 32'd4997;
    weight_rom[45][52] = 32'd3216;
    weight_rom[45][53] = -32'd1245;
    weight_rom[45][54] = 32'd2323;
    weight_rom[45][55] = -32'd6312;
    weight_rom[45][56] = 32'd119;
    weight_rom[45][57] = -32'd1359;
    weight_rom[45][58] = -32'd2173;
    weight_rom[45][59] = -32'd6399;
    weight_rom[45][60] = -32'd4722;
    weight_rom[45][61] = -32'd2677;
    weight_rom[45][62] = -32'd3787;
    weight_rom[45][63] = 32'd3544;
    weight_rom[46][0] = -32'd2467;
    weight_rom[46][1] = 32'd1902;
    weight_rom[46][2] = 32'd532;
    weight_rom[46][3] = -32'd4679;
    weight_rom[46][4] = 32'd3344;
    weight_rom[46][5] = 32'd938;
    weight_rom[46][6] = 32'd4848;
    weight_rom[46][7] = 32'd1984;
    weight_rom[46][8] = -32'd2669;
    weight_rom[46][9] = 32'd3272;
    weight_rom[46][10] = -32'd4166;
    weight_rom[46][11] = -32'd6155;
    weight_rom[46][12] = 32'd1238;
    weight_rom[46][13] = -32'd4560;
    weight_rom[46][14] = 32'd5610;
    weight_rom[46][15] = -32'd4135;
    weight_rom[46][16] = -32'd2789;
    weight_rom[46][17] = -32'd5288;
    weight_rom[46][18] = 32'd1783;
    weight_rom[46][19] = -32'd4917;
    weight_rom[46][20] = -32'd5939;
    weight_rom[46][21] = 32'd5802;
    weight_rom[46][22] = 32'd5904;
    weight_rom[46][23] = -32'd4204;
    weight_rom[46][24] = -32'd3298;
    weight_rom[46][25] = 32'd1;
    weight_rom[46][26] = 32'd4127;
    weight_rom[46][27] = 32'd6517;
    weight_rom[46][28] = 32'd3280;
    weight_rom[46][29] = -32'd918;
    weight_rom[46][30] = 32'd5458;
    weight_rom[46][31] = 32'd1854;
    weight_rom[46][32] = -32'd5316;
    weight_rom[46][33] = 32'd1949;
    weight_rom[46][34] = -32'd4326;
    weight_rom[46][35] = 32'd3274;
    weight_rom[46][36] = -32'd1528;
    weight_rom[46][37] = 32'd728;
    weight_rom[46][38] = 32'd5039;
    weight_rom[46][39] = 32'd2983;
    weight_rom[46][40] = -32'd3812;
    weight_rom[46][41] = 32'd3597;
    weight_rom[46][42] = 32'd6224;
    weight_rom[46][43] = -32'd3145;
    weight_rom[46][44] = 32'd2781;
    weight_rom[46][45] = -32'd2067;
    weight_rom[46][46] = -32'd1449;
    weight_rom[46][47] = -32'd105;
    weight_rom[46][48] = 32'd2587;
    weight_rom[46][49] = 32'd1936;
    weight_rom[46][50] = 32'd6144;
    weight_rom[46][51] = -32'd5532;
    weight_rom[46][52] = -32'd1586;
    weight_rom[46][53] = 32'd5656;
    weight_rom[46][54] = 32'd2655;
    weight_rom[46][55] = 32'd2018;
    weight_rom[46][56] = -32'd4620;
    weight_rom[46][57] = 32'd2541;
    weight_rom[46][58] = 32'd4166;
    weight_rom[46][59] = 32'd6519;
    weight_rom[46][60] = -32'd5293;
    weight_rom[46][61] = -32'd56;
    weight_rom[46][62] = 32'd2468;
    weight_rom[46][63] = -32'd4;
    weight_rom[47][0] = 32'd263;
    weight_rom[47][1] = -32'd4268;
    weight_rom[47][2] = 32'd1801;
    weight_rom[47][3] = 32'd3427;
    weight_rom[47][4] = 32'd1576;
    weight_rom[47][5] = -32'd2883;
    weight_rom[47][6] = 32'd246;
    weight_rom[47][7] = 32'd4321;
    weight_rom[47][8] = -32'd3491;
    weight_rom[47][9] = -32'd4848;
    weight_rom[47][10] = 32'd3797;
    weight_rom[47][11] = 32'd5648;
    weight_rom[47][12] = -32'd42;
    weight_rom[47][13] = -32'd5749;
    weight_rom[47][14] = -32'd3609;
    weight_rom[47][15] = -32'd1805;
    weight_rom[47][16] = 32'd3838;
    weight_rom[47][17] = -32'd3383;
    weight_rom[47][18] = 32'd5417;
    weight_rom[47][19] = 32'd3856;
    weight_rom[47][20] = -32'd2933;
    weight_rom[47][21] = 32'd3738;
    weight_rom[47][22] = 32'd1069;
    weight_rom[47][23] = 32'd3932;
    weight_rom[47][24] = -32'd3743;
    weight_rom[47][25] = -32'd1153;
    weight_rom[47][26] = 32'd3644;
    weight_rom[47][27] = -32'd6160;
    weight_rom[47][28] = -32'd4560;
    weight_rom[47][29] = 32'd4337;
    weight_rom[47][30] = 32'd1774;
    weight_rom[47][31] = -32'd3147;
    weight_rom[47][32] = 32'd4345;
    weight_rom[47][33] = 32'd5958;
    weight_rom[47][34] = -32'd4889;
    weight_rom[47][35] = 32'd5413;
    weight_rom[47][36] = -32'd4347;
    weight_rom[47][37] = -32'd2734;
    weight_rom[47][38] = 32'd707;
    weight_rom[47][39] = 32'd5539;
    weight_rom[47][40] = -32'd4845;
    weight_rom[47][41] = -32'd4791;
    weight_rom[47][42] = -32'd1165;
    weight_rom[47][43] = -32'd1506;
    weight_rom[47][44] = -32'd4248;
    weight_rom[47][45] = 32'd6309;
    weight_rom[47][46] = 32'd3048;
    weight_rom[47][47] = 32'd953;
    weight_rom[47][48] = 32'd1871;
    weight_rom[47][49] = -32'd6169;
    weight_rom[47][50] = -32'd206;
    weight_rom[47][51] = 32'd2710;
    weight_rom[47][52] = -32'd2585;
    weight_rom[47][53] = -32'd5386;
    weight_rom[47][54] = 32'd5976;
    weight_rom[47][55] = 32'd1554;
    weight_rom[47][56] = 32'd1463;
    weight_rom[47][57] = -32'd139;
    weight_rom[47][58] = -32'd6050;
    weight_rom[47][59] = -32'd2869;
    weight_rom[47][60] = -32'd988;
    weight_rom[47][61] = -32'd1033;
    weight_rom[47][62] = -32'd3673;
    weight_rom[47][63] = -32'd2553;
    weight_rom[48][0] = 32'd612;
    weight_rom[48][1] = 32'd2502;
    weight_rom[48][2] = 32'd2963;
    weight_rom[48][3] = 32'd1549;
    weight_rom[48][4] = 32'd2674;
    weight_rom[48][5] = 32'd3532;
    weight_rom[48][6] = 32'd1196;
    weight_rom[48][7] = -32'd3848;
    weight_rom[48][8] = -32'd6001;
    weight_rom[48][9] = 32'd3385;
    weight_rom[48][10] = 32'd2080;
    weight_rom[48][11] = 32'd2484;
    weight_rom[48][12] = 32'd6393;
    weight_rom[48][13] = 32'd3679;
    weight_rom[48][14] = -32'd1675;
    weight_rom[48][15] = -32'd2169;
    weight_rom[48][16] = 32'd1017;
    weight_rom[48][17] = -32'd6391;
    weight_rom[48][18] = 32'd1475;
    weight_rom[48][19] = -32'd2939;
    weight_rom[48][20] = 32'd2712;
    weight_rom[48][21] = 32'd6439;
    weight_rom[48][22] = -32'd830;
    weight_rom[48][23] = 32'd690;
    weight_rom[48][24] = -32'd3004;
    weight_rom[48][25] = 32'd4856;
    weight_rom[48][26] = 32'd3419;
    weight_rom[48][27] = 32'd5208;
    weight_rom[48][28] = -32'd546;
    weight_rom[48][29] = -32'd4982;
    weight_rom[48][30] = 32'd1701;
    weight_rom[48][31] = 32'd5060;
    weight_rom[48][32] = 32'd5484;
    weight_rom[48][33] = -32'd4568;
    weight_rom[48][34] = -32'd4937;
    weight_rom[48][35] = 32'd945;
    weight_rom[48][36] = 32'd4409;
    weight_rom[48][37] = -32'd1082;
    weight_rom[48][38] = 32'd452;
    weight_rom[48][39] = 32'd3436;
    weight_rom[48][40] = -32'd3885;
    weight_rom[48][41] = -32'd423;
    weight_rom[48][42] = -32'd724;
    weight_rom[48][43] = 32'd5806;
    weight_rom[48][44] = -32'd3468;
    weight_rom[48][45] = 32'd1699;
    weight_rom[48][46] = 32'd2421;
    weight_rom[48][47] = -32'd3429;
    weight_rom[48][48] = 32'd3705;
    weight_rom[48][49] = 32'd1548;
    weight_rom[48][50] = -32'd5719;
    weight_rom[48][51] = 32'd5505;
    weight_rom[48][52] = -32'd532;
    weight_rom[48][53] = 32'd151;
    weight_rom[48][54] = 32'd410;
    weight_rom[48][55] = -32'd2492;
    weight_rom[48][56] = 32'd861;
    weight_rom[48][57] = 32'd164;
    weight_rom[48][58] = 32'd4860;
    weight_rom[48][59] = 32'd2202;
    weight_rom[48][60] = 32'd5684;
    weight_rom[48][61] = -32'd1172;
    weight_rom[48][62] = -32'd803;
    weight_rom[48][63] = 32'd6209;
    weight_rom[49][0] = -32'd4130;
    weight_rom[49][1] = -32'd1484;
    weight_rom[49][2] = 32'd6237;
    weight_rom[49][3] = -32'd5228;
    weight_rom[49][4] = -32'd3762;
    weight_rom[49][5] = -32'd4101;
    weight_rom[49][6] = -32'd1323;
    weight_rom[49][7] = -32'd6409;
    weight_rom[49][8] = -32'd6319;
    weight_rom[49][9] = -32'd6231;
    weight_rom[49][10] = -32'd23;
    weight_rom[49][11] = 32'd2313;
    weight_rom[49][12] = -32'd4765;
    weight_rom[49][13] = -32'd526;
    weight_rom[49][14] = -32'd890;
    weight_rom[49][15] = -32'd6210;
    weight_rom[49][16] = 32'd1763;
    weight_rom[49][17] = -32'd409;
    weight_rom[49][18] = 32'd4898;
    weight_rom[49][19] = 32'd4942;
    weight_rom[49][20] = -32'd5731;
    weight_rom[49][21] = 32'd583;
    weight_rom[49][22] = 32'd1049;
    weight_rom[49][23] = -32'd1355;
    weight_rom[49][24] = -32'd3308;
    weight_rom[49][25] = 32'd1722;
    weight_rom[49][26] = -32'd4093;
    weight_rom[49][27] = 32'd1607;
    weight_rom[49][28] = -32'd1950;
    weight_rom[49][29] = 32'd3079;
    weight_rom[49][30] = -32'd1268;
    weight_rom[49][31] = 32'd5186;
    weight_rom[49][32] = 32'd1963;
    weight_rom[49][33] = -32'd296;
    weight_rom[49][34] = 32'd243;
    weight_rom[49][35] = -32'd4184;
    weight_rom[49][36] = 32'd641;
    weight_rom[49][37] = -32'd1613;
    weight_rom[49][38] = -32'd3991;
    weight_rom[49][39] = 32'd1202;
    weight_rom[49][40] = 32'd3526;
    weight_rom[49][41] = 32'd1387;
    weight_rom[49][42] = 32'd1003;
    weight_rom[49][43] = 32'd1446;
    weight_rom[49][44] = -32'd73;
    weight_rom[49][45] = -32'd1098;
    weight_rom[49][46] = -32'd3773;
    weight_rom[49][47] = 32'd3852;
    weight_rom[49][48] = 32'd5734;
    weight_rom[49][49] = 32'd124;
    weight_rom[49][50] = 32'd677;
    weight_rom[49][51] = -32'd3005;
    weight_rom[49][52] = 32'd4167;
    weight_rom[49][53] = 32'd5485;
    weight_rom[49][54] = -32'd1314;
    weight_rom[49][55] = -32'd5429;
    weight_rom[49][56] = 32'd2814;
    weight_rom[49][57] = -32'd3043;
    weight_rom[49][58] = 32'd167;
    weight_rom[49][59] = -32'd4237;
    weight_rom[49][60] = 32'd555;
    weight_rom[49][61] = -32'd3521;
    weight_rom[49][62] = 32'd3696;
    weight_rom[49][63] = 32'd2141;
    weight_rom[50][0] = 32'd6154;
    weight_rom[50][1] = 32'd5724;
    weight_rom[50][2] = 32'd213;
    weight_rom[50][3] = -32'd5451;
    weight_rom[50][4] = -32'd4766;
    weight_rom[50][5] = -32'd2311;
    weight_rom[50][6] = -32'd5835;
    weight_rom[50][7] = -32'd4759;
    weight_rom[50][8] = 32'd6392;
    weight_rom[50][9] = -32'd6263;
    weight_rom[50][10] = 32'd725;
    weight_rom[50][11] = -32'd3726;
    weight_rom[50][12] = 32'd2557;
    weight_rom[50][13] = -32'd5791;
    weight_rom[50][14] = -32'd794;
    weight_rom[50][15] = -32'd6236;
    weight_rom[50][16] = 32'd3904;
    weight_rom[50][17] = -32'd2604;
    weight_rom[50][18] = 32'd2935;
    weight_rom[50][19] = 32'd5820;
    weight_rom[50][20] = 32'd4447;
    weight_rom[50][21] = 32'd6065;
    weight_rom[50][22] = 32'd218;
    weight_rom[50][23] = -32'd4827;
    weight_rom[50][24] = -32'd5734;
    weight_rom[50][25] = 32'd426;
    weight_rom[50][26] = -32'd5395;
    weight_rom[50][27] = 32'd6204;
    weight_rom[50][28] = -32'd5324;
    weight_rom[50][29] = 32'd412;
    weight_rom[50][30] = 32'd3308;
    weight_rom[50][31] = -32'd2657;
    weight_rom[50][32] = -32'd5197;
    weight_rom[50][33] = 32'd1334;
    weight_rom[50][34] = -32'd3331;
    weight_rom[50][35] = -32'd3030;
    weight_rom[50][36] = -32'd4073;
    weight_rom[50][37] = 32'd4927;
    weight_rom[50][38] = -32'd4374;
    weight_rom[50][39] = -32'd4036;
    weight_rom[50][40] = -32'd976;
    weight_rom[50][41] = -32'd939;
    weight_rom[50][42] = 32'd6335;
    weight_rom[50][43] = 32'd4390;
    weight_rom[50][44] = 32'd5437;
    weight_rom[50][45] = -32'd4370;
    weight_rom[50][46] = -32'd3420;
    weight_rom[50][47] = -32'd177;
    weight_rom[50][48] = 32'd2515;
    weight_rom[50][49] = 32'd599;
    weight_rom[50][50] = 32'd4470;
    weight_rom[50][51] = -32'd1697;
    weight_rom[50][52] = 32'd5635;
    weight_rom[50][53] = 32'd5296;
    weight_rom[50][54] = 32'd5946;
    weight_rom[50][55] = -32'd5361;
    weight_rom[50][56] = 32'd5737;
    weight_rom[50][57] = -32'd590;
    weight_rom[50][58] = -32'd1333;
    weight_rom[50][59] = 32'd1051;
    weight_rom[50][60] = 32'd359;
    weight_rom[50][61] = -32'd4766;
    weight_rom[50][62] = 32'd3721;
    weight_rom[50][63] = -32'd1202;
    weight_rom[51][0] = 32'd3606;
    weight_rom[51][1] = -32'd4751;
    weight_rom[51][2] = -32'd2320;
    weight_rom[51][3] = 32'd2634;
    weight_rom[51][4] = -32'd6362;
    weight_rom[51][5] = -32'd977;
    weight_rom[51][6] = -32'd2160;
    weight_rom[51][7] = 32'd5243;
    weight_rom[51][8] = -32'd946;
    weight_rom[51][9] = -32'd2311;
    weight_rom[51][10] = 32'd2873;
    weight_rom[51][11] = 32'd2082;
    weight_rom[51][12] = -32'd1254;
    weight_rom[51][13] = 32'd6486;
    weight_rom[51][14] = 32'd1480;
    weight_rom[51][15] = 32'd4347;
    weight_rom[51][16] = -32'd1363;
    weight_rom[51][17] = 32'd1289;
    weight_rom[51][18] = -32'd4973;
    weight_rom[51][19] = -32'd4603;
    weight_rom[51][20] = -32'd6503;
    weight_rom[51][21] = -32'd5562;
    weight_rom[51][22] = 32'd3391;
    weight_rom[51][23] = 32'd4787;
    weight_rom[51][24] = -32'd538;
    weight_rom[51][25] = -32'd5041;
    weight_rom[51][26] = 32'd2607;
    weight_rom[51][27] = -32'd458;
    weight_rom[51][28] = -32'd181;
    weight_rom[51][29] = -32'd2779;
    weight_rom[51][30] = 32'd410;
    weight_rom[51][31] = -32'd3539;
    weight_rom[51][32] = -32'd1284;
    weight_rom[51][33] = 32'd1071;
    weight_rom[51][34] = -32'd1859;
    weight_rom[51][35] = -32'd3949;
    weight_rom[51][36] = 32'd2888;
    weight_rom[51][37] = 32'd5312;
    weight_rom[51][38] = 32'd5459;
    weight_rom[51][39] = 32'd2184;
    weight_rom[51][40] = 32'd857;
    weight_rom[51][41] = -32'd6198;
    weight_rom[51][42] = -32'd3386;
    weight_rom[51][43] = 32'd2757;
    weight_rom[51][44] = -32'd3778;
    weight_rom[51][45] = 32'd6372;
    weight_rom[51][46] = -32'd2866;
    weight_rom[51][47] = -32'd2175;
    weight_rom[51][48] = -32'd4510;
    weight_rom[51][49] = -32'd1842;
    weight_rom[51][50] = 32'd6512;
    weight_rom[51][51] = 32'd903;
    weight_rom[51][52] = 32'd590;
    weight_rom[51][53] = -32'd4501;
    weight_rom[51][54] = 32'd1862;
    weight_rom[51][55] = 32'd5547;
    weight_rom[51][56] = 32'd5403;
    weight_rom[51][57] = -32'd382;
    weight_rom[51][58] = -32'd37;
    weight_rom[51][59] = 32'd5295;
    weight_rom[51][60] = -32'd4703;
    weight_rom[51][61] = -32'd3975;
    weight_rom[51][62] = -32'd612;
    weight_rom[51][63] = -32'd2877;
    weight_rom[52][0] = 32'd5760;
    weight_rom[52][1] = -32'd2083;
    weight_rom[52][2] = 32'd3869;
    weight_rom[52][3] = -32'd5599;
    weight_rom[52][4] = -32'd1958;
    weight_rom[52][5] = 32'd99;
    weight_rom[52][6] = 32'd3969;
    weight_rom[52][7] = 32'd4900;
    weight_rom[52][8] = -32'd1516;
    weight_rom[52][9] = -32'd148;
    weight_rom[52][10] = -32'd3559;
    weight_rom[52][11] = -32'd1391;
    weight_rom[52][12] = -32'd941;
    weight_rom[52][13] = -32'd5796;
    weight_rom[52][14] = 32'd5807;
    weight_rom[52][15] = -32'd2974;
    weight_rom[52][16] = 32'd5440;
    weight_rom[52][17] = -32'd2657;
    weight_rom[52][18] = 32'd5275;
    weight_rom[52][19] = -32'd489;
    weight_rom[52][20] = -32'd3318;
    weight_rom[52][21] = -32'd1760;
    weight_rom[52][22] = -32'd2850;
    weight_rom[52][23] = -32'd4492;
    weight_rom[52][24] = 32'd3050;
    weight_rom[52][25] = 32'd1384;
    weight_rom[52][26] = -32'd1725;
    weight_rom[52][27] = 32'd4553;
    weight_rom[52][28] = 32'd5514;
    weight_rom[52][29] = -32'd94;
    weight_rom[52][30] = 32'd2325;
    weight_rom[52][31] = -32'd1162;
    weight_rom[52][32] = 32'd3000;
    weight_rom[52][33] = -32'd1291;
    weight_rom[52][34] = 32'd6416;
    weight_rom[52][35] = -32'd3318;
    weight_rom[52][36] = 32'd145;
    weight_rom[52][37] = -32'd92;
    weight_rom[52][38] = -32'd2256;
    weight_rom[52][39] = 32'd1617;
    weight_rom[52][40] = -32'd6278;
    weight_rom[52][41] = 32'd3715;
    weight_rom[52][42] = 32'd2376;
    weight_rom[52][43] = -32'd5078;
    weight_rom[52][44] = -32'd4663;
    weight_rom[52][45] = 32'd4205;
    weight_rom[52][46] = -32'd1164;
    weight_rom[52][47] = -32'd5153;
    weight_rom[52][48] = -32'd3362;
    weight_rom[52][49] = -32'd5485;
    weight_rom[52][50] = -32'd912;
    weight_rom[52][51] = 32'd5003;
    weight_rom[52][52] = 32'd2116;
    weight_rom[52][53] = -32'd1747;
    weight_rom[52][54] = -32'd2645;
    weight_rom[52][55] = 32'd2480;
    weight_rom[52][56] = 32'd5846;
    weight_rom[52][57] = 32'd2708;
    weight_rom[52][58] = 32'd2194;
    weight_rom[52][59] = -32'd2356;
    weight_rom[52][60] = -32'd6543;
    weight_rom[52][61] = -32'd5828;
    weight_rom[52][62] = 32'd3829;
    weight_rom[52][63] = 32'd3029;
    weight_rom[53][0] = 32'd5175;
    weight_rom[53][1] = -32'd5066;
    weight_rom[53][2] = -32'd3003;
    weight_rom[53][3] = 32'd4218;
    weight_rom[53][4] = 32'd1178;
    weight_rom[53][5] = -32'd3376;
    weight_rom[53][6] = -32'd6492;
    weight_rom[53][7] = 32'd1276;
    weight_rom[53][8] = 32'd2354;
    weight_rom[53][9] = 32'd3544;
    weight_rom[53][10] = 32'd6505;
    weight_rom[53][11] = 32'd1982;
    weight_rom[53][12] = 32'd2852;
    weight_rom[53][13] = 32'd2556;
    weight_rom[53][14] = -32'd3398;
    weight_rom[53][15] = 32'd236;
    weight_rom[53][16] = 32'd432;
    weight_rom[53][17] = -32'd2622;
    weight_rom[53][18] = -32'd5682;
    weight_rom[53][19] = 32'd6304;
    weight_rom[53][20] = 32'd3157;
    weight_rom[53][21] = -32'd3599;
    weight_rom[53][22] = -32'd1926;
    weight_rom[53][23] = -32'd2493;
    weight_rom[53][24] = 32'd1398;
    weight_rom[53][25] = -32'd5017;
    weight_rom[53][26] = -32'd886;
    weight_rom[53][27] = -32'd5735;
    weight_rom[53][28] = -32'd6028;
    weight_rom[53][29] = -32'd2622;
    weight_rom[53][30] = -32'd937;
    weight_rom[53][31] = -32'd3400;
    weight_rom[53][32] = 32'd3667;
    weight_rom[53][33] = -32'd2122;
    weight_rom[53][34] = 32'd2415;
    weight_rom[53][35] = -32'd2537;
    weight_rom[53][36] = 32'd1367;
    weight_rom[53][37] = -32'd2226;
    weight_rom[53][38] = -32'd1676;
    weight_rom[53][39] = 32'd1343;
    weight_rom[53][40] = -32'd6102;
    weight_rom[53][41] = -32'd6415;
    weight_rom[53][42] = 32'd2830;
    weight_rom[53][43] = 32'd3092;
    weight_rom[53][44] = 32'd3394;
    weight_rom[53][45] = -32'd2864;
    weight_rom[53][46] = -32'd3482;
    weight_rom[53][47] = -32'd3423;
    weight_rom[53][48] = 32'd4485;
    weight_rom[53][49] = -32'd4019;
    weight_rom[53][50] = -32'd2355;
    weight_rom[53][51] = 32'd5792;
    weight_rom[53][52] = 32'd5285;
    weight_rom[53][53] = 32'd1561;
    weight_rom[53][54] = -32'd4895;
    weight_rom[53][55] = -32'd4887;
    weight_rom[53][56] = -32'd3346;
    weight_rom[53][57] = 32'd5775;
    weight_rom[53][58] = -32'd6386;
    weight_rom[53][59] = 32'd2231;
    weight_rom[53][60] = 32'd4065;
    weight_rom[53][61] = -32'd3956;
    weight_rom[53][62] = 32'd4438;
    weight_rom[53][63] = -32'd3379;
    weight_rom[54][0] = 32'd1283;
    weight_rom[54][1] = 32'd5566;
    weight_rom[54][2] = -32'd799;
    weight_rom[54][3] = 32'd2703;
    weight_rom[54][4] = -32'd1412;
    weight_rom[54][5] = -32'd5048;
    weight_rom[54][6] = -32'd2182;
    weight_rom[54][7] = 32'd1317;
    weight_rom[54][8] = -32'd3692;
    weight_rom[54][9] = 32'd2402;
    weight_rom[54][10] = 32'd6223;
    weight_rom[54][11] = -32'd5156;
    weight_rom[54][12] = 32'd2522;
    weight_rom[54][13] = 32'd6339;
    weight_rom[54][14] = -32'd4961;
    weight_rom[54][15] = -32'd2638;
    weight_rom[54][16] = -32'd4483;
    weight_rom[54][17] = 32'd3187;
    weight_rom[54][18] = 32'd445;
    weight_rom[54][19] = -32'd217;
    weight_rom[54][20] = -32'd2408;
    weight_rom[54][21] = -32'd3986;
    weight_rom[54][22] = 32'd5165;
    weight_rom[54][23] = -32'd2751;
    weight_rom[54][24] = 32'd2265;
    weight_rom[54][25] = -32'd2133;
    weight_rom[54][26] = -32'd6145;
    weight_rom[54][27] = -32'd2159;
    weight_rom[54][28] = -32'd2733;
    weight_rom[54][29] = 32'd1259;
    weight_rom[54][30] = 32'd3034;
    weight_rom[54][31] = 32'd2259;
    weight_rom[54][32] = -32'd5004;
    weight_rom[54][33] = -32'd4891;
    weight_rom[54][34] = 32'd5884;
    weight_rom[54][35] = 32'd722;
    weight_rom[54][36] = -32'd512;
    weight_rom[54][37] = -32'd5153;
    weight_rom[54][38] = 32'd3405;
    weight_rom[54][39] = -32'd133;
    weight_rom[54][40] = -32'd710;
    weight_rom[54][41] = 32'd3432;
    weight_rom[54][42] = 32'd1406;
    weight_rom[54][43] = -32'd2947;
    weight_rom[54][44] = 32'd8;
    weight_rom[54][45] = -32'd5635;
    weight_rom[54][46] = -32'd6296;
    weight_rom[54][47] = 32'd5888;
    weight_rom[54][48] = -32'd3810;
    weight_rom[54][49] = 32'd5908;
    weight_rom[54][50] = 32'd5330;
    weight_rom[54][51] = 32'd3140;
    weight_rom[54][52] = -32'd5261;
    weight_rom[54][53] = -32'd4464;
    weight_rom[54][54] = 32'd4489;
    weight_rom[54][55] = -32'd1877;
    weight_rom[54][56] = -32'd4829;
    weight_rom[54][57] = -32'd2237;
    weight_rom[54][58] = 32'd4869;
    weight_rom[54][59] = -32'd4090;
    weight_rom[54][60] = -32'd5405;
    weight_rom[54][61] = -32'd6433;
    weight_rom[54][62] = 32'd2028;
    weight_rom[54][63] = -32'd4302;
    weight_rom[55][0] = 32'd5529;
    weight_rom[55][1] = 32'd4945;
    weight_rom[55][2] = -32'd5525;
    weight_rom[55][3] = -32'd5487;
    weight_rom[55][4] = -32'd819;
    weight_rom[55][5] = 32'd1449;
    weight_rom[55][6] = -32'd1334;
    weight_rom[55][7] = 32'd2163;
    weight_rom[55][8] = 32'd5897;
    weight_rom[55][9] = -32'd709;
    weight_rom[55][10] = 32'd1970;
    weight_rom[55][11] = 32'd2068;
    weight_rom[55][12] = 32'd6438;
    weight_rom[55][13] = -32'd3418;
    weight_rom[55][14] = -32'd3965;
    weight_rom[55][15] = 32'd5776;
    weight_rom[55][16] = 32'd2567;
    weight_rom[55][17] = -32'd5922;
    weight_rom[55][18] = -32'd4690;
    weight_rom[55][19] = 32'd4765;
    weight_rom[55][20] = -32'd5218;
    weight_rom[55][21] = -32'd4708;
    weight_rom[55][22] = 32'd5851;
    weight_rom[55][23] = 32'd4868;
    weight_rom[55][24] = -32'd5489;
    weight_rom[55][25] = -32'd4681;
    weight_rom[55][26] = -32'd3151;
    weight_rom[55][27] = -32'd5675;
    weight_rom[55][28] = -32'd3833;
    weight_rom[55][29] = -32'd867;
    weight_rom[55][30] = 32'd4252;
    weight_rom[55][31] = 32'd4273;
    weight_rom[55][32] = -32'd6553;
    weight_rom[55][33] = -32'd1418;
    weight_rom[55][34] = -32'd4685;
    weight_rom[55][35] = 32'd1153;
    weight_rom[55][36] = 32'd4308;
    weight_rom[55][37] = 32'd5942;
    weight_rom[55][38] = -32'd2112;
    weight_rom[55][39] = 32'd375;
    weight_rom[55][40] = 32'd4150;
    weight_rom[55][41] = 32'd5155;
    weight_rom[55][42] = -32'd5392;
    weight_rom[55][43] = 32'd1823;
    weight_rom[55][44] = 32'd5397;
    weight_rom[55][45] = -32'd5811;
    weight_rom[55][46] = 32'd4972;
    weight_rom[55][47] = -32'd2554;
    weight_rom[55][48] = -32'd5603;
    weight_rom[55][49] = -32'd1196;
    weight_rom[55][50] = -32'd4046;
    weight_rom[55][51] = -32'd5418;
    weight_rom[55][52] = -32'd3511;
    weight_rom[55][53] = 32'd6134;
    weight_rom[55][54] = -32'd1806;
    weight_rom[55][55] = 32'd1212;
    weight_rom[55][56] = -32'd2591;
    weight_rom[55][57] = -32'd6000;
    weight_rom[55][58] = -32'd698;
    weight_rom[55][59] = 32'd1635;
    weight_rom[55][60] = 32'd1754;
    weight_rom[55][61] = 32'd1668;
    weight_rom[55][62] = -32'd3559;
    weight_rom[55][63] = 32'd391;
    weight_rom[56][0] = -32'd5393;
    weight_rom[56][1] = -32'd3172;
    weight_rom[56][2] = -32'd6221;
    weight_rom[56][3] = -32'd5441;
    weight_rom[56][4] = 32'd5297;
    weight_rom[56][5] = -32'd2770;
    weight_rom[56][6] = 32'd490;
    weight_rom[56][7] = -32'd4254;
    weight_rom[56][8] = 32'd3753;
    weight_rom[56][9] = -32'd2967;
    weight_rom[56][10] = -32'd3938;
    weight_rom[56][11] = 32'd6545;
    weight_rom[56][12] = -32'd4870;
    weight_rom[56][13] = -32'd4689;
    weight_rom[56][14] = 32'd5071;
    weight_rom[56][15] = -32'd3154;
    weight_rom[56][16] = 32'd3843;
    weight_rom[56][17] = 32'd5280;
    weight_rom[56][18] = -32'd6400;
    weight_rom[56][19] = 32'd1163;
    weight_rom[56][20] = -32'd1831;
    weight_rom[56][21] = 32'd1604;
    weight_rom[56][22] = 32'd5145;
    weight_rom[56][23] = 32'd2263;
    weight_rom[56][24] = 32'd5917;
    weight_rom[56][25] = 32'd2517;
    weight_rom[56][26] = -32'd6112;
    weight_rom[56][27] = 32'd6230;
    weight_rom[56][28] = -32'd3432;
    weight_rom[56][29] = -32'd4398;
    weight_rom[56][30] = -32'd4634;
    weight_rom[56][31] = 32'd2268;
    weight_rom[56][32] = 32'd2780;
    weight_rom[56][33] = -32'd4421;
    weight_rom[56][34] = -32'd1544;
    weight_rom[56][35] = -32'd963;
    weight_rom[56][36] = 32'd4319;
    weight_rom[56][37] = -32'd5764;
    weight_rom[56][38] = 32'd5925;
    weight_rom[56][39] = -32'd2169;
    weight_rom[56][40] = 32'd5049;
    weight_rom[56][41] = -32'd880;
    weight_rom[56][42] = 32'd2318;
    weight_rom[56][43] = -32'd2084;
    weight_rom[56][44] = -32'd4631;
    weight_rom[56][45] = -32'd4975;
    weight_rom[56][46] = 32'd6102;
    weight_rom[56][47] = -32'd4340;
    weight_rom[56][48] = 32'd2664;
    weight_rom[56][49] = -32'd436;
    weight_rom[56][50] = 32'd1512;
    weight_rom[56][51] = 32'd2217;
    weight_rom[56][52] = 32'd2738;
    weight_rom[56][53] = 32'd5436;
    weight_rom[56][54] = 32'd2103;
    weight_rom[56][55] = 32'd4398;
    weight_rom[56][56] = 32'd5178;
    weight_rom[56][57] = -32'd48;
    weight_rom[56][58] = -32'd2058;
    weight_rom[56][59] = -32'd2143;
    weight_rom[56][60] = 32'd5434;
    weight_rom[56][61] = -32'd2406;
    weight_rom[56][62] = -32'd2962;
    weight_rom[56][63] = -32'd2752;
    weight_rom[57][0] = -32'd3984;
    weight_rom[57][1] = 32'd2096;
    weight_rom[57][2] = 32'd6064;
    weight_rom[57][3] = 32'd6378;
    weight_rom[57][4] = -32'd1988;
    weight_rom[57][5] = 32'd1064;
    weight_rom[57][6] = 32'd5503;
    weight_rom[57][7] = 32'd5431;
    weight_rom[57][8] = -32'd5381;
    weight_rom[57][9] = 32'd6515;
    weight_rom[57][10] = 32'd2362;
    weight_rom[57][11] = -32'd5921;
    weight_rom[57][12] = -32'd5189;
    weight_rom[57][13] = -32'd4962;
    weight_rom[57][14] = 32'd1911;
    weight_rom[57][15] = -32'd922;
    weight_rom[57][16] = -32'd2401;
    weight_rom[57][17] = 32'd4617;
    weight_rom[57][18] = -32'd1021;
    weight_rom[57][19] = -32'd1634;
    weight_rom[57][20] = -32'd3009;
    weight_rom[57][21] = 32'd3687;
    weight_rom[57][22] = -32'd1055;
    weight_rom[57][23] = 32'd3888;
    weight_rom[57][24] = 32'd4436;
    weight_rom[57][25] = -32'd3850;
    weight_rom[57][26] = 32'd4970;
    weight_rom[57][27] = 32'd4154;
    weight_rom[57][28] = 32'd5353;
    weight_rom[57][29] = -32'd5025;
    weight_rom[57][30] = 32'd4363;
    weight_rom[57][31] = 32'd4251;
    weight_rom[57][32] = -32'd1879;
    weight_rom[57][33] = 32'd3071;
    weight_rom[57][34] = 32'd717;
    weight_rom[57][35] = 32'd1512;
    weight_rom[57][36] = 32'd2744;
    weight_rom[57][37] = -32'd2652;
    weight_rom[57][38] = 32'd3118;
    weight_rom[57][39] = 32'd253;
    weight_rom[57][40] = -32'd5417;
    weight_rom[57][41] = 32'd465;
    weight_rom[57][42] = -32'd5713;
    weight_rom[57][43] = 32'd6523;
    weight_rom[57][44] = 32'd1912;
    weight_rom[57][45] = 32'd1058;
    weight_rom[57][46] = -32'd2076;
    weight_rom[57][47] = -32'd515;
    weight_rom[57][48] = -32'd1277;
    weight_rom[57][49] = -32'd5862;
    weight_rom[57][50] = -32'd1235;
    weight_rom[57][51] = -32'd1175;
    weight_rom[57][52] = 32'd4243;
    weight_rom[57][53] = -32'd4365;
    weight_rom[57][54] = -32'd382;
    weight_rom[57][55] = -32'd5981;
    weight_rom[57][56] = 32'd6187;
    weight_rom[57][57] = 32'd582;
    weight_rom[57][58] = -32'd4741;
    weight_rom[57][59] = -32'd3785;
    weight_rom[57][60] = -32'd3818;
    weight_rom[57][61] = 32'd6201;
    weight_rom[57][62] = -32'd2426;
    weight_rom[57][63] = 32'd1689;
    weight_rom[58][0] = -32'd5960;
    weight_rom[58][1] = 32'd4157;
    weight_rom[58][2] = 32'd4403;
    weight_rom[58][3] = -32'd1647;
    weight_rom[58][4] = 32'd183;
    weight_rom[58][5] = -32'd4530;
    weight_rom[58][6] = -32'd2013;
    weight_rom[58][7] = -32'd1064;
    weight_rom[58][8] = -32'd1080;
    weight_rom[58][9] = -32'd967;
    weight_rom[58][10] = -32'd5607;
    weight_rom[58][11] = 32'd6254;
    weight_rom[58][12] = 32'd2940;
    weight_rom[58][13] = -32'd2578;
    weight_rom[58][14] = -32'd2806;
    weight_rom[58][15] = 32'd4885;
    weight_rom[58][16] = 32'd4681;
    weight_rom[58][17] = 32'd2199;
    weight_rom[58][18] = -32'd2686;
    weight_rom[58][19] = -32'd2807;
    weight_rom[58][20] = 32'd4491;
    weight_rom[58][21] = 32'd1026;
    weight_rom[58][22] = 32'd3674;
    weight_rom[58][23] = -32'd3270;
    weight_rom[58][24] = 32'd3998;
    weight_rom[58][25] = -32'd1417;
    weight_rom[58][26] = -32'd3363;
    weight_rom[58][27] = 32'd4620;
    weight_rom[58][28] = -32'd418;
    weight_rom[58][29] = 32'd612;
    weight_rom[58][30] = 32'd528;
    weight_rom[58][31] = -32'd1350;
    weight_rom[58][32] = -32'd3218;
    weight_rom[58][33] = -32'd3816;
    weight_rom[58][34] = -32'd5547;
    weight_rom[58][35] = -32'd5484;
    weight_rom[58][36] = -32'd5172;
    weight_rom[58][37] = -32'd2646;
    weight_rom[58][38] = 32'd1277;
    weight_rom[58][39] = -32'd3964;
    weight_rom[58][40] = 32'd502;
    weight_rom[58][41] = -32'd301;
    weight_rom[58][42] = 32'd1260;
    weight_rom[58][43] = -32'd3099;
    weight_rom[58][44] = -32'd3501;
    weight_rom[58][45] = 32'd5619;
    weight_rom[58][46] = -32'd2116;
    weight_rom[58][47] = -32'd2528;
    weight_rom[58][48] = 32'd5505;
    weight_rom[58][49] = -32'd6061;
    weight_rom[58][50] = -32'd6015;
    weight_rom[58][51] = -32'd384;
    weight_rom[58][52] = 32'd4679;
    weight_rom[58][53] = -32'd4965;
    weight_rom[58][54] = -32'd3946;
    weight_rom[58][55] = -32'd3451;
    weight_rom[58][56] = 32'd4709;
    weight_rom[58][57] = -32'd4345;
    weight_rom[58][58] = -32'd793;
    weight_rom[58][59] = -32'd2448;
    weight_rom[58][60] = 32'd2166;
    weight_rom[58][61] = -32'd4014;
    weight_rom[58][62] = -32'd5022;
    weight_rom[58][63] = -32'd5007;
    weight_rom[59][0] = -32'd2289;
    weight_rom[59][1] = 32'd723;
    weight_rom[59][2] = 32'd2568;
    weight_rom[59][3] = -32'd1695;
    weight_rom[59][4] = 32'd3717;
    weight_rom[59][5] = -32'd247;
    weight_rom[59][6] = -32'd2005;
    weight_rom[59][7] = -32'd1531;
    weight_rom[59][8] = 32'd4969;
    weight_rom[59][9] = -32'd637;
    weight_rom[59][10] = -32'd6151;
    weight_rom[59][11] = -32'd1220;
    weight_rom[59][12] = 32'd1027;
    weight_rom[59][13] = -32'd5229;
    weight_rom[59][14] = 32'd4141;
    weight_rom[59][15] = 32'd4481;
    weight_rom[59][16] = 32'd5323;
    weight_rom[59][17] = 32'd1221;
    weight_rom[59][18] = -32'd183;
    weight_rom[59][19] = -32'd3889;
    weight_rom[59][20] = -32'd2446;
    weight_rom[59][21] = -32'd4627;
    weight_rom[59][22] = -32'd310;
    weight_rom[59][23] = 32'd1636;
    weight_rom[59][24] = 32'd4233;
    weight_rom[59][25] = 32'd5186;
    weight_rom[59][26] = 32'd751;
    weight_rom[59][27] = 32'd5740;
    weight_rom[59][28] = -32'd441;
    weight_rom[59][29] = 32'd5274;
    weight_rom[59][30] = 32'd4517;
    weight_rom[59][31] = -32'd4504;
    weight_rom[59][32] = -32'd6384;
    weight_rom[59][33] = -32'd5785;
    weight_rom[59][34] = -32'd6498;
    weight_rom[59][35] = -32'd5402;
    weight_rom[59][36] = 32'd4441;
    weight_rom[59][37] = -32'd2354;
    weight_rom[59][38] = 32'd4992;
    weight_rom[59][39] = 32'd3999;
    weight_rom[59][40] = 32'd5416;
    weight_rom[59][41] = -32'd1452;
    weight_rom[59][42] = 32'd3140;
    weight_rom[59][43] = -32'd2894;
    weight_rom[59][44] = -32'd4498;
    weight_rom[59][45] = -32'd42;
    weight_rom[59][46] = -32'd6460;
    weight_rom[59][47] = -32'd6092;
    weight_rom[59][48] = 32'd1969;
    weight_rom[59][49] = 32'd2846;
    weight_rom[59][50] = -32'd2001;
    weight_rom[59][51] = -32'd5909;
    weight_rom[59][52] = -32'd1112;
    weight_rom[59][53] = -32'd5434;
    weight_rom[59][54] = 32'd1332;
    weight_rom[59][55] = 32'd5108;
    weight_rom[59][56] = -32'd5111;
    weight_rom[59][57] = 32'd3413;
    weight_rom[59][58] = -32'd48;
    weight_rom[59][59] = -32'd4209;
    weight_rom[59][60] = -32'd5522;
    weight_rom[59][61] = -32'd2020;
    weight_rom[59][62] = -32'd2973;
    weight_rom[59][63] = 32'd2030;
    weight_rom[60][0] = -32'd1459;
    weight_rom[60][1] = 32'd388;
    weight_rom[60][2] = -32'd1193;
    weight_rom[60][3] = 32'd4099;
    weight_rom[60][4] = -32'd1356;
    weight_rom[60][5] = 32'd427;
    weight_rom[60][6] = 32'd3112;
    weight_rom[60][7] = 32'd247;
    weight_rom[60][8] = 32'd5829;
    weight_rom[60][9] = -32'd4408;
    weight_rom[60][10] = -32'd3176;
    weight_rom[60][11] = 32'd4859;
    weight_rom[60][12] = -32'd2960;
    weight_rom[60][13] = 32'd2518;
    weight_rom[60][14] = 32'd4736;
    weight_rom[60][15] = -32'd4114;
    weight_rom[60][16] = -32'd2924;
    weight_rom[60][17] = 32'd5141;
    weight_rom[60][18] = 32'd1011;
    weight_rom[60][19] = 32'd3431;
    weight_rom[60][20] = 32'd3787;
    weight_rom[60][21] = 32'd4077;
    weight_rom[60][22] = -32'd32;
    weight_rom[60][23] = 32'd940;
    weight_rom[60][24] = 32'd5671;
    weight_rom[60][25] = -32'd3875;
    weight_rom[60][26] = -32'd6042;
    weight_rom[60][27] = -32'd5438;
    weight_rom[60][28] = 32'd3415;
    weight_rom[60][29] = -32'd2045;
    weight_rom[60][30] = -32'd900;
    weight_rom[60][31] = 32'd3118;
    weight_rom[60][32] = 32'd528;
    weight_rom[60][33] = 32'd686;
    weight_rom[60][34] = 32'd2233;
    weight_rom[60][35] = -32'd4301;
    weight_rom[60][36] = 32'd2241;
    weight_rom[60][37] = -32'd4400;
    weight_rom[60][38] = -32'd5903;
    weight_rom[60][39] = -32'd4118;
    weight_rom[60][40] = -32'd1468;
    weight_rom[60][41] = 32'd5078;
    weight_rom[60][42] = -32'd3788;
    weight_rom[60][43] = 32'd5644;
    weight_rom[60][44] = 32'd2404;
    weight_rom[60][45] = 32'd4495;
    weight_rom[60][46] = 32'd2362;
    weight_rom[60][47] = -32'd2318;
    weight_rom[60][48] = -32'd5368;
    weight_rom[60][49] = 32'd499;
    weight_rom[60][50] = -32'd3077;
    weight_rom[60][51] = -32'd4049;
    weight_rom[60][52] = -32'd5382;
    weight_rom[60][53] = 32'd5366;
    weight_rom[60][54] = -32'd5758;
    weight_rom[60][55] = -32'd6433;
    weight_rom[60][56] = 32'd5864;
    weight_rom[60][57] = 32'd6356;
    weight_rom[60][58] = -32'd1262;
    weight_rom[60][59] = 32'd5267;
    weight_rom[60][60] = 32'd1359;
    weight_rom[60][61] = -32'd1863;
    weight_rom[60][62] = -32'd3807;
    weight_rom[60][63] = -32'd2840;
    weight_rom[61][0] = -32'd2996;
    weight_rom[61][1] = -32'd3383;
    weight_rom[61][2] = -32'd4282;
    weight_rom[61][3] = 32'd5862;
    weight_rom[61][4] = 32'd1600;
    weight_rom[61][5] = -32'd5874;
    weight_rom[61][6] = -32'd626;
    weight_rom[61][7] = -32'd5938;
    weight_rom[61][8] = -32'd427;
    weight_rom[61][9] = 32'd3864;
    weight_rom[61][10] = -32'd489;
    weight_rom[61][11] = 32'd3701;
    weight_rom[61][12] = -32'd5512;
    weight_rom[61][13] = -32'd5737;
    weight_rom[61][14] = 32'd4541;
    weight_rom[61][15] = 32'd3966;
    weight_rom[61][16] = 32'd6337;
    weight_rom[61][17] = -32'd4124;
    weight_rom[61][18] = -32'd5980;
    weight_rom[61][19] = -32'd1487;
    weight_rom[61][20] = 32'd5136;
    weight_rom[61][21] = 32'd1781;
    weight_rom[61][22] = -32'd3870;
    weight_rom[61][23] = 32'd4362;
    weight_rom[61][24] = 32'd580;
    weight_rom[61][25] = 32'd102;
    weight_rom[61][26] = 32'd2186;
    weight_rom[61][27] = -32'd1499;
    weight_rom[61][28] = -32'd4528;
    weight_rom[61][29] = 32'd3053;
    weight_rom[61][30] = -32'd1585;
    weight_rom[61][31] = -32'd1828;
    weight_rom[61][32] = 32'd4602;
    weight_rom[61][33] = 32'd1248;
    weight_rom[61][34] = 32'd1858;
    weight_rom[61][35] = 32'd236;
    weight_rom[61][36] = 32'd2582;
    weight_rom[61][37] = 32'd3711;
    weight_rom[61][38] = -32'd3184;
    weight_rom[61][39] = -32'd5439;
    weight_rom[61][40] = 32'd4319;
    weight_rom[61][41] = 32'd5163;
    weight_rom[61][42] = 32'd4477;
    weight_rom[61][43] = -32'd6230;
    weight_rom[61][44] = 32'd1227;
    weight_rom[61][45] = -32'd709;
    weight_rom[61][46] = 32'd4265;
    weight_rom[61][47] = 32'd578;
    weight_rom[61][48] = 32'd5870;
    weight_rom[61][49] = 32'd114;
    weight_rom[61][50] = 32'd2439;
    weight_rom[61][51] = 32'd3807;
    weight_rom[61][52] = -32'd815;
    weight_rom[61][53] = -32'd4015;
    weight_rom[61][54] = -32'd1135;
    weight_rom[61][55] = -32'd3913;
    weight_rom[61][56] = -32'd1004;
    weight_rom[61][57] = 32'd5842;
    weight_rom[61][58] = 32'd2341;
    weight_rom[61][59] = -32'd1347;
    weight_rom[61][60] = -32'd4404;
    weight_rom[61][61] = -32'd6442;
    weight_rom[61][62] = -32'd585;
    weight_rom[61][63] = -32'd6550;
    weight_rom[62][0] = 32'd4308;
    weight_rom[62][1] = -32'd5333;
    weight_rom[62][2] = -32'd4503;
    weight_rom[62][3] = 32'd6370;
    weight_rom[62][4] = 32'd4749;
    weight_rom[62][5] = -32'd2141;
    weight_rom[62][6] = -32'd3609;
    weight_rom[62][7] = -32'd4374;
    weight_rom[62][8] = 32'd1486;
    weight_rom[62][9] = 32'd2538;
    weight_rom[62][10] = 32'd4827;
    weight_rom[62][11] = 32'd878;
    weight_rom[62][12] = -32'd5430;
    weight_rom[62][13] = 32'd123;
    weight_rom[62][14] = 32'd5490;
    weight_rom[62][15] = -32'd548;
    weight_rom[62][16] = -32'd4709;
    weight_rom[62][17] = -32'd5518;
    weight_rom[62][18] = -32'd4941;
    weight_rom[62][19] = 32'd147;
    weight_rom[62][20] = -32'd867;
    weight_rom[62][21] = -32'd1465;
    weight_rom[62][22] = 32'd1194;
    weight_rom[62][23] = 32'd5322;
    weight_rom[62][24] = -32'd3928;
    weight_rom[62][25] = -32'd1058;
    weight_rom[62][26] = -32'd2319;
    weight_rom[62][27] = -32'd5622;
    weight_rom[62][28] = -32'd166;
    weight_rom[62][29] = 32'd2079;
    weight_rom[62][30] = 32'd5440;
    weight_rom[62][31] = 32'd2244;
    weight_rom[62][32] = 32'd5998;
    weight_rom[62][33] = 32'd4874;
    weight_rom[62][34] = -32'd1169;
    weight_rom[62][35] = -32'd3748;
    weight_rom[62][36] = -32'd1795;
    weight_rom[62][37] = -32'd4947;
    weight_rom[62][38] = -32'd458;
    weight_rom[62][39] = -32'd835;
    weight_rom[62][40] = -32'd4801;
    weight_rom[62][41] = -32'd2152;
    weight_rom[62][42] = -32'd6155;
    weight_rom[62][43] = 32'd2578;
    weight_rom[62][44] = 32'd3340;
    weight_rom[62][45] = 32'd2733;
    weight_rom[62][46] = -32'd4631;
    weight_rom[62][47] = 32'd677;
    weight_rom[62][48] = -32'd3164;
    weight_rom[62][49] = -32'd3366;
    weight_rom[62][50] = 32'd5882;
    weight_rom[62][51] = -32'd603;
    weight_rom[62][52] = -32'd3529;
    weight_rom[62][53] = -32'd1097;
    weight_rom[62][54] = 32'd610;
    weight_rom[62][55] = 32'd6016;
    weight_rom[62][56] = -32'd6431;
    weight_rom[62][57] = -32'd3970;
    weight_rom[62][58] = -32'd1036;
    weight_rom[62][59] = -32'd3338;
    weight_rom[62][60] = 32'd3092;
    weight_rom[62][61] = 32'd4446;
    weight_rom[62][62] = 32'd5353;
    weight_rom[62][63] = -32'd4889;
    weight_rom[63][0] = -32'd1877;
    weight_rom[63][1] = 32'd5206;
    weight_rom[63][2] = -32'd3273;
    weight_rom[63][3] = 32'd3321;
    weight_rom[63][4] = 32'd5891;
    weight_rom[63][5] = -32'd4791;
    weight_rom[63][6] = -32'd623;
    weight_rom[63][7] = 32'd3119;
    weight_rom[63][8] = -32'd4364;
    weight_rom[63][9] = -32'd3659;
    weight_rom[63][10] = 32'd2977;
    weight_rom[63][11] = 32'd3125;
    weight_rom[63][12] = 32'd5166;
    weight_rom[63][13] = 32'd6510;
    weight_rom[63][14] = -32'd3247;
    weight_rom[63][15] = -32'd223;
    weight_rom[63][16] = -32'd3905;
    weight_rom[63][17] = -32'd3414;
    weight_rom[63][18] = 32'd768;
    weight_rom[63][19] = -32'd100;
    weight_rom[63][20] = 32'd5373;
    weight_rom[63][21] = 32'd2282;
    weight_rom[63][22] = -32'd4113;
    weight_rom[63][23] = -32'd6394;
    weight_rom[63][24] = 32'd1530;
    weight_rom[63][25] = -32'd6316;
    weight_rom[63][26] = 32'd5215;
    weight_rom[63][27] = -32'd3790;
    weight_rom[63][28] = -32'd917;
    weight_rom[63][29] = 32'd5656;
    weight_rom[63][30] = -32'd3261;
    weight_rom[63][31] = -32'd3006;
    weight_rom[63][32] = 32'd861;
    weight_rom[63][33] = 32'd1008;
    weight_rom[63][34] = -32'd135;
    weight_rom[63][35] = -32'd2840;
    weight_rom[63][36] = 32'd4971;
    weight_rom[63][37] = 32'd1768;
    weight_rom[63][38] = -32'd3578;
    weight_rom[63][39] = 32'd2074;
    weight_rom[63][40] = 32'd5706;
    weight_rom[63][41] = 32'd1508;
    weight_rom[63][42] = 32'd4506;
    weight_rom[63][43] = 32'd2953;
    weight_rom[63][44] = -32'd2497;
    weight_rom[63][45] = 32'd3039;
    weight_rom[63][46] = -32'd4460;
    weight_rom[63][47] = -32'd1880;
    weight_rom[63][48] = -32'd2133;
    weight_rom[63][49] = 32'd3207;
    weight_rom[63][50] = -32'd3040;
    weight_rom[63][51] = -32'd2599;
    weight_rom[63][52] = -32'd2736;
    weight_rom[63][53] = -32'd670;
    weight_rom[63][54] = -32'd838;
    weight_rom[63][55] = 32'd1486;
    weight_rom[63][56] = -32'd755;
    weight_rom[63][57] = 32'd4919;
    weight_rom[63][58] = 32'd6047;
    weight_rom[63][59] = -32'd676;
    weight_rom[63][60] = -32'd2605;
    weight_rom[63][61] = -32'd6134;
    weight_rom[63][62] = -32'd5184;
    weight_rom[63][63] = 32'd5683;
    weight_rom[64][0] = -32'd2871;
    weight_rom[64][1] = 32'd5248;
    weight_rom[64][2] = 32'd645;
    weight_rom[64][3] = -32'd1621;
    weight_rom[64][4] = -32'd4625;
    weight_rom[64][5] = -32'd5722;
    weight_rom[64][6] = -32'd4707;
    weight_rom[64][7] = -32'd5468;
    weight_rom[64][8] = 32'd6437;
    weight_rom[64][9] = -32'd5473;
    weight_rom[64][10] = 32'd3181;
    weight_rom[64][11] = 32'd4961;
    weight_rom[64][12] = -32'd4038;
    weight_rom[64][13] = 32'd4115;
    weight_rom[64][14] = 32'd3342;
    weight_rom[64][15] = -32'd4804;
    weight_rom[64][16] = -32'd4138;
    weight_rom[64][17] = 32'd3861;
    weight_rom[64][18] = -32'd2055;
    weight_rom[64][19] = 32'd1012;
    weight_rom[64][20] = -32'd1607;
    weight_rom[64][21] = -32'd3146;
    weight_rom[64][22] = -32'd2207;
    weight_rom[64][23] = 32'd2280;
    weight_rom[64][24] = 32'd3183;
    weight_rom[64][25] = 32'd3837;
    weight_rom[64][26] = 32'd5087;
    weight_rom[64][27] = -32'd3547;
    weight_rom[64][28] = 32'd1270;
    weight_rom[64][29] = 32'd4207;
    weight_rom[64][30] = 32'd4511;
    weight_rom[64][31] = -32'd5488;
    weight_rom[64][32] = 32'd189;
    weight_rom[64][33] = -32'd2025;
    weight_rom[64][34] = -32'd1108;
    weight_rom[64][35] = -32'd1306;
    weight_rom[64][36] = 32'd2953;
    weight_rom[64][37] = -32'd4930;
    weight_rom[64][38] = 32'd3196;
    weight_rom[64][39] = -32'd816;
    weight_rom[64][40] = 32'd3295;
    weight_rom[64][41] = 32'd5595;
    weight_rom[64][42] = -32'd519;
    weight_rom[64][43] = 32'd4409;
    weight_rom[64][44] = -32'd681;
    weight_rom[64][45] = -32'd4273;
    weight_rom[64][46] = 32'd3802;
    weight_rom[64][47] = -32'd690;
    weight_rom[64][48] = -32'd1281;
    weight_rom[64][49] = -32'd4348;
    weight_rom[64][50] = 32'd4082;
    weight_rom[64][51] = -32'd1520;
    weight_rom[64][52] = 32'd3568;
    weight_rom[64][53] = 32'd1297;
    weight_rom[64][54] = 32'd3259;
    weight_rom[64][55] = -32'd3123;
    weight_rom[64][56] = -32'd5949;
    weight_rom[64][57] = 32'd2680;
    weight_rom[64][58] = 32'd1301;
    weight_rom[64][59] = -32'd2352;
    weight_rom[64][60] = -32'd479;
    weight_rom[64][61] = 32'd5769;
    weight_rom[64][62] = 32'd2887;
    weight_rom[64][63] = 32'd4814;
    weight_rom[65][0] = 32'd559;
    weight_rom[65][1] = 32'd1744;
    weight_rom[65][2] = 32'd2812;
    weight_rom[65][3] = -32'd5459;
    weight_rom[65][4] = 32'd5591;
    weight_rom[65][5] = 32'd6422;
    weight_rom[65][6] = -32'd4241;
    weight_rom[65][7] = 32'd1352;
    weight_rom[65][8] = -32'd3517;
    weight_rom[65][9] = 32'd2365;
    weight_rom[65][10] = -32'd976;
    weight_rom[65][11] = -32'd1256;
    weight_rom[65][12] = -32'd2315;
    weight_rom[65][13] = 32'd1510;
    weight_rom[65][14] = -32'd517;
    weight_rom[65][15] = -32'd5497;
    weight_rom[65][16] = 32'd5164;
    weight_rom[65][17] = -32'd6099;
    weight_rom[65][18] = 32'd3003;
    weight_rom[65][19] = 32'd4791;
    weight_rom[65][20] = 32'd6082;
    weight_rom[65][21] = -32'd2029;
    weight_rom[65][22] = 32'd4653;
    weight_rom[65][23] = -32'd5874;
    weight_rom[65][24] = 32'd3118;
    weight_rom[65][25] = -32'd5648;
    weight_rom[65][26] = -32'd2289;
    weight_rom[65][27] = -32'd404;
    weight_rom[65][28] = 32'd6547;
    weight_rom[65][29] = 32'd873;
    weight_rom[65][30] = -32'd209;
    weight_rom[65][31] = 32'd6456;
    weight_rom[65][32] = -32'd5438;
    weight_rom[65][33] = 32'd3971;
    weight_rom[65][34] = -32'd6238;
    weight_rom[65][35] = 32'd4087;
    weight_rom[65][36] = -32'd5077;
    weight_rom[65][37] = -32'd5629;
    weight_rom[65][38] = 32'd5494;
    weight_rom[65][39] = -32'd2926;
    weight_rom[65][40] = 32'd5784;
    weight_rom[65][41] = 32'd6056;
    weight_rom[65][42] = -32'd3701;
    weight_rom[65][43] = 32'd6218;
    weight_rom[65][44] = -32'd1239;
    weight_rom[65][45] = -32'd1819;
    weight_rom[65][46] = 32'd1524;
    weight_rom[65][47] = 32'd6101;
    weight_rom[65][48] = -32'd5882;
    weight_rom[65][49] = -32'd4064;
    weight_rom[65][50] = -32'd5827;
    weight_rom[65][51] = 32'd4645;
    weight_rom[65][52] = -32'd5563;
    weight_rom[65][53] = -32'd5613;
    weight_rom[65][54] = 32'd4298;
    weight_rom[65][55] = -32'd5675;
    weight_rom[65][56] = 32'd575;
    weight_rom[65][57] = -32'd604;
    weight_rom[65][58] = 32'd4030;
    weight_rom[65][59] = 32'd3203;
    weight_rom[65][60] = 32'd1303;
    weight_rom[65][61] = 32'd5139;
    weight_rom[65][62] = 32'd2454;
    weight_rom[65][63] = -32'd3491;
    weight_rom[66][0] = -32'd4706;
    weight_rom[66][1] = -32'd2109;
    weight_rom[66][2] = 32'd2099;
    weight_rom[66][3] = 32'd3632;
    weight_rom[66][4] = -32'd103;
    weight_rom[66][5] = -32'd2328;
    weight_rom[66][6] = -32'd21;
    weight_rom[66][7] = -32'd3337;
    weight_rom[66][8] = 32'd5802;
    weight_rom[66][9] = 32'd2025;
    weight_rom[66][10] = -32'd2019;
    weight_rom[66][11] = -32'd2267;
    weight_rom[66][12] = -32'd3582;
    weight_rom[66][13] = -32'd2539;
    weight_rom[66][14] = 32'd4482;
    weight_rom[66][15] = 32'd2987;
    weight_rom[66][16] = 32'd2022;
    weight_rom[66][17] = 32'd1085;
    weight_rom[66][18] = 32'd1996;
    weight_rom[66][19] = 32'd6301;
    weight_rom[66][20] = -32'd5383;
    weight_rom[66][21] = 32'd5472;
    weight_rom[66][22] = -32'd3839;
    weight_rom[66][23] = 32'd640;
    weight_rom[66][24] = 32'd281;
    weight_rom[66][25] = -32'd337;
    weight_rom[66][26] = 32'd5255;
    weight_rom[66][27] = -32'd3033;
    weight_rom[66][28] = 32'd3531;
    weight_rom[66][29] = 32'd2058;
    weight_rom[66][30] = 32'd184;
    weight_rom[66][31] = -32'd4506;
    weight_rom[66][32] = 32'd640;
    weight_rom[66][33] = 32'd527;
    weight_rom[66][34] = -32'd2157;
    weight_rom[66][35] = -32'd6371;
    weight_rom[66][36] = -32'd1208;
    weight_rom[66][37] = 32'd5366;
    weight_rom[66][38] = -32'd999;
    weight_rom[66][39] = 32'd762;
    weight_rom[66][40] = 32'd2314;
    weight_rom[66][41] = 32'd117;
    weight_rom[66][42] = -32'd4800;
    weight_rom[66][43] = 32'd6233;
    weight_rom[66][44] = 32'd6345;
    weight_rom[66][45] = 32'd1799;
    weight_rom[66][46] = -32'd5965;
    weight_rom[66][47] = -32'd1607;
    weight_rom[66][48] = -32'd45;
    weight_rom[66][49] = -32'd514;
    weight_rom[66][50] = 32'd499;
    weight_rom[66][51] = 32'd3263;
    weight_rom[66][52] = 32'd4293;
    weight_rom[66][53] = -32'd3581;
    weight_rom[66][54] = 32'd3555;
    weight_rom[66][55] = -32'd6184;
    weight_rom[66][56] = -32'd2116;
    weight_rom[66][57] = 32'd532;
    weight_rom[66][58] = -32'd5120;
    weight_rom[66][59] = 32'd6176;
    weight_rom[66][60] = -32'd4308;
    weight_rom[66][61] = 32'd465;
    weight_rom[66][62] = -32'd5298;
    weight_rom[66][63] = 32'd3648;
    weight_rom[67][0] = 32'd3960;
    weight_rom[67][1] = -32'd1976;
    weight_rom[67][2] = -32'd2884;
    weight_rom[67][3] = 32'd765;
    weight_rom[67][4] = -32'd3168;
    weight_rom[67][5] = 32'd4061;
    weight_rom[67][6] = -32'd1062;
    weight_rom[67][7] = -32'd1451;
    weight_rom[67][8] = 32'd1961;
    weight_rom[67][9] = -32'd2971;
    weight_rom[67][10] = -32'd1690;
    weight_rom[67][11] = 32'd2196;
    weight_rom[67][12] = -32'd1900;
    weight_rom[67][13] = 32'd1623;
    weight_rom[67][14] = 32'd2994;
    weight_rom[67][15] = -32'd46;
    weight_rom[67][16] = -32'd4559;
    weight_rom[67][17] = 32'd6493;
    weight_rom[67][18] = 32'd4529;
    weight_rom[67][19] = -32'd1211;
    weight_rom[67][20] = 32'd2451;
    weight_rom[67][21] = -32'd2745;
    weight_rom[67][22] = -32'd5620;
    weight_rom[67][23] = -32'd2783;
    weight_rom[67][24] = -32'd5656;
    weight_rom[67][25] = 32'd795;
    weight_rom[67][26] = 32'd6503;
    weight_rom[67][27] = -32'd5230;
    weight_rom[67][28] = -32'd1338;
    weight_rom[67][29] = 32'd5221;
    weight_rom[67][30] = -32'd2510;
    weight_rom[67][31] = 32'd6401;
    weight_rom[67][32] = -32'd1573;
    weight_rom[67][33] = -32'd5514;
    weight_rom[67][34] = -32'd4232;
    weight_rom[67][35] = 32'd1957;
    weight_rom[67][36] = 32'd5064;
    weight_rom[67][37] = -32'd4061;
    weight_rom[67][38] = -32'd2069;
    weight_rom[67][39] = -32'd2005;
    weight_rom[67][40] = -32'd1790;
    weight_rom[67][41] = -32'd618;
    weight_rom[67][42] = 32'd5941;
    weight_rom[67][43] = -32'd5698;
    weight_rom[67][44] = -32'd2723;
    weight_rom[67][45] = -32'd5626;
    weight_rom[67][46] = 32'd1606;
    weight_rom[67][47] = -32'd3168;
    weight_rom[67][48] = -32'd4937;
    weight_rom[67][49] = -32'd2801;
    weight_rom[67][50] = -32'd5628;
    weight_rom[67][51] = -32'd2984;
    weight_rom[67][52] = -32'd948;
    weight_rom[67][53] = 32'd5655;
    weight_rom[67][54] = -32'd6044;
    weight_rom[67][55] = -32'd3345;
    weight_rom[67][56] = -32'd348;
    weight_rom[67][57] = 32'd4582;
    weight_rom[67][58] = -32'd1346;
    weight_rom[67][59] = -32'd812;
    weight_rom[67][60] = 32'd3167;
    weight_rom[67][61] = 32'd571;
    weight_rom[67][62] = 32'd5538;
    weight_rom[67][63] = 32'd1423;
    weight_rom[68][0] = -32'd5576;
    weight_rom[68][1] = 32'd2961;
    weight_rom[68][2] = 32'd5962;
    weight_rom[68][3] = -32'd993;
    weight_rom[68][4] = -32'd535;
    weight_rom[68][5] = -32'd3215;
    weight_rom[68][6] = 32'd5437;
    weight_rom[68][7] = -32'd2769;
    weight_rom[68][8] = 32'd1412;
    weight_rom[68][9] = 32'd5909;
    weight_rom[68][10] = 32'd6391;
    weight_rom[68][11] = 32'd4034;
    weight_rom[68][12] = -32'd5643;
    weight_rom[68][13] = 32'd354;
    weight_rom[68][14] = 32'd3623;
    weight_rom[68][15] = -32'd827;
    weight_rom[68][16] = -32'd782;
    weight_rom[68][17] = 32'd4662;
    weight_rom[68][18] = 32'd2523;
    weight_rom[68][19] = 32'd4292;
    weight_rom[68][20] = -32'd81;
    weight_rom[68][21] = -32'd393;
    weight_rom[68][22] = -32'd5649;
    weight_rom[68][23] = -32'd2532;
    weight_rom[68][24] = -32'd1689;
    weight_rom[68][25] = 32'd1683;
    weight_rom[68][26] = 32'd4265;
    weight_rom[68][27] = -32'd4358;
    weight_rom[68][28] = 32'd4293;
    weight_rom[68][29] = -32'd1317;
    weight_rom[68][30] = 32'd957;
    weight_rom[68][31] = 32'd6255;
    weight_rom[68][32] = 32'd1404;
    weight_rom[68][33] = 32'd863;
    weight_rom[68][34] = -32'd5263;
    weight_rom[68][35] = 32'd2213;
    weight_rom[68][36] = -32'd5935;
    weight_rom[68][37] = 32'd4210;
    weight_rom[68][38] = 32'd6049;
    weight_rom[68][39] = 32'd5673;
    weight_rom[68][40] = 32'd5743;
    weight_rom[68][41] = -32'd2900;
    weight_rom[68][42] = -32'd5601;
    weight_rom[68][43] = 32'd4218;
    weight_rom[68][44] = -32'd2689;
    weight_rom[68][45] = -32'd1814;
    weight_rom[68][46] = -32'd2504;
    weight_rom[68][47] = -32'd3362;
    weight_rom[68][48] = -32'd1298;
    weight_rom[68][49] = -32'd3310;
    weight_rom[68][50] = 32'd5688;
    weight_rom[68][51] = -32'd5013;
    weight_rom[68][52] = 32'd1259;
    weight_rom[68][53] = 32'd5353;
    weight_rom[68][54] = -32'd4009;
    weight_rom[68][55] = 32'd5000;
    weight_rom[68][56] = 32'd1483;
    weight_rom[68][57] = -32'd260;
    weight_rom[68][58] = -32'd2138;
    weight_rom[68][59] = 32'd4732;
    weight_rom[68][60] = -32'd2586;
    weight_rom[68][61] = 32'd2015;
    weight_rom[68][62] = 32'd897;
    weight_rom[68][63] = 32'd6172;
    weight_rom[69][0] = 32'd6381;
    weight_rom[69][1] = 32'd5205;
    weight_rom[69][2] = 32'd3118;
    weight_rom[69][3] = 32'd5326;
    weight_rom[69][4] = 32'd6291;
    weight_rom[69][5] = 32'd2379;
    weight_rom[69][6] = -32'd1803;
    weight_rom[69][7] = -32'd1891;
    weight_rom[69][8] = 32'd166;
    weight_rom[69][9] = -32'd4573;
    weight_rom[69][10] = -32'd6027;
    weight_rom[69][11] = 32'd3437;
    weight_rom[69][12] = 32'd249;
    weight_rom[69][13] = -32'd968;
    weight_rom[69][14] = 32'd2046;
    weight_rom[69][15] = 32'd3008;
    weight_rom[69][16] = 32'd1511;
    weight_rom[69][17] = 32'd281;
    weight_rom[69][18] = -32'd918;
    weight_rom[69][19] = 32'd3467;
    weight_rom[69][20] = -32'd1472;
    weight_rom[69][21] = 32'd5113;
    weight_rom[69][22] = 32'd5777;
    weight_rom[69][23] = -32'd1927;
    weight_rom[69][24] = 32'd5515;
    weight_rom[69][25] = 32'd2472;
    weight_rom[69][26] = 32'd4520;
    weight_rom[69][27] = -32'd4623;
    weight_rom[69][28] = -32'd4316;
    weight_rom[69][29] = -32'd2270;
    weight_rom[69][30] = -32'd2291;
    weight_rom[69][31] = 32'd3851;
    weight_rom[69][32] = -32'd1458;
    weight_rom[69][33] = 32'd5347;
    weight_rom[69][34] = 32'd5986;
    weight_rom[69][35] = 32'd3914;
    weight_rom[69][36] = 32'd6047;
    weight_rom[69][37] = 32'd584;
    weight_rom[69][38] = -32'd722;
    weight_rom[69][39] = 32'd5539;
    weight_rom[69][40] = -32'd2941;
    weight_rom[69][41] = 32'd6014;
    weight_rom[69][42] = -32'd3944;
    weight_rom[69][43] = 32'd1917;
    weight_rom[69][44] = -32'd1906;
    weight_rom[69][45] = 32'd456;
    weight_rom[69][46] = -32'd1720;
    weight_rom[69][47] = -32'd553;
    weight_rom[69][48] = -32'd1956;
    weight_rom[69][49] = 32'd1903;
    weight_rom[69][50] = 32'd3491;
    weight_rom[69][51] = -32'd3250;
    weight_rom[69][52] = -32'd5378;
    weight_rom[69][53] = 32'd3686;
    weight_rom[69][54] = 32'd479;
    weight_rom[69][55] = -32'd1102;
    weight_rom[69][56] = 32'd4833;
    weight_rom[69][57] = -32'd1661;
    weight_rom[69][58] = 32'd910;
    weight_rom[69][59] = 32'd863;
    weight_rom[69][60] = 32'd2128;
    weight_rom[69][61] = -32'd1480;
    weight_rom[69][62] = -32'd1786;
    weight_rom[69][63] = -32'd1656;
    weight_rom[70][0] = 32'd3568;
    weight_rom[70][1] = 32'd5073;
    weight_rom[70][2] = 32'd712;
    weight_rom[70][3] = -32'd5096;
    weight_rom[70][4] = -32'd96;
    weight_rom[70][5] = 32'd3410;
    weight_rom[70][6] = 32'd1056;
    weight_rom[70][7] = 32'd2871;
    weight_rom[70][8] = -32'd3530;
    weight_rom[70][9] = -32'd886;
    weight_rom[70][10] = 32'd4810;
    weight_rom[70][11] = 32'd3903;
    weight_rom[70][12] = -32'd5667;
    weight_rom[70][13] = -32'd4840;
    weight_rom[70][14] = -32'd4227;
    weight_rom[70][15] = 32'd3480;
    weight_rom[70][16] = -32'd5459;
    weight_rom[70][17] = -32'd5719;
    weight_rom[70][18] = 32'd2267;
    weight_rom[70][19] = 32'd963;
    weight_rom[70][20] = 32'd1739;
    weight_rom[70][21] = 32'd2722;
    weight_rom[70][22] = 32'd90;
    weight_rom[70][23] = 32'd1589;
    weight_rom[70][24] = 32'd1106;
    weight_rom[70][25] = -32'd3233;
    weight_rom[70][26] = -32'd3289;
    weight_rom[70][27] = 32'd6200;
    weight_rom[70][28] = -32'd6154;
    weight_rom[70][29] = -32'd6411;
    weight_rom[70][30] = -32'd6038;
    weight_rom[70][31] = 32'd2089;
    weight_rom[70][32] = -32'd3403;
    weight_rom[70][33] = -32'd1359;
    weight_rom[70][34] = 32'd1302;
    weight_rom[70][35] = 32'd5672;
    weight_rom[70][36] = 32'd2348;
    weight_rom[70][37] = -32'd5533;
    weight_rom[70][38] = -32'd143;
    weight_rom[70][39] = 32'd31;
    weight_rom[70][40] = -32'd2199;
    weight_rom[70][41] = -32'd4681;
    weight_rom[70][42] = -32'd1994;
    weight_rom[70][43] = 32'd1931;
    weight_rom[70][44] = 32'd846;
    weight_rom[70][45] = 32'd6504;
    weight_rom[70][46] = 32'd3535;
    weight_rom[70][47] = 32'd3401;
    weight_rom[70][48] = 32'd3576;
    weight_rom[70][49] = 32'd1978;
    weight_rom[70][50] = 32'd2070;
    weight_rom[70][51] = 32'd5514;
    weight_rom[70][52] = -32'd2131;
    weight_rom[70][53] = -32'd6299;
    weight_rom[70][54] = 32'd5699;
    weight_rom[70][55] = 32'd2887;
    weight_rom[70][56] = 32'd2122;
    weight_rom[70][57] = -32'd88;
    weight_rom[70][58] = 32'd4733;
    weight_rom[70][59] = -32'd4492;
    weight_rom[70][60] = -32'd4478;
    weight_rom[70][61] = 32'd1929;
    weight_rom[70][62] = 32'd3362;
    weight_rom[70][63] = 32'd2378;
    weight_rom[71][0] = -32'd3949;
    weight_rom[71][1] = 32'd3668;
    weight_rom[71][2] = 32'd1464;
    weight_rom[71][3] = -32'd96;
    weight_rom[71][4] = -32'd2244;
    weight_rom[71][5] = 32'd1253;
    weight_rom[71][6] = 32'd1733;
    weight_rom[71][7] = -32'd2659;
    weight_rom[71][8] = -32'd4239;
    weight_rom[71][9] = 32'd5814;
    weight_rom[71][10] = 32'd1031;
    weight_rom[71][11] = -32'd844;
    weight_rom[71][12] = 32'd3936;
    weight_rom[71][13] = 32'd5067;
    weight_rom[71][14] = 32'd590;
    weight_rom[71][15] = -32'd4470;
    weight_rom[71][16] = 32'd5012;
    weight_rom[71][17] = 32'd4343;
    weight_rom[71][18] = -32'd2944;
    weight_rom[71][19] = 32'd5977;
    weight_rom[71][20] = 32'd2671;
    weight_rom[71][21] = -32'd5738;
    weight_rom[71][22] = -32'd1187;
    weight_rom[71][23] = -32'd2175;
    weight_rom[71][24] = 32'd502;
    weight_rom[71][25] = -32'd6422;
    weight_rom[71][26] = 32'd1005;
    weight_rom[71][27] = 32'd3398;
    weight_rom[71][28] = -32'd3873;
    weight_rom[71][29] = 32'd4280;
    weight_rom[71][30] = -32'd2988;
    weight_rom[71][31] = 32'd1019;
    weight_rom[71][32] = -32'd5308;
    weight_rom[71][33] = -32'd2669;
    weight_rom[71][34] = 32'd2997;
    weight_rom[71][35] = -32'd6289;
    weight_rom[71][36] = 32'd1721;
    weight_rom[71][37] = 32'd5969;
    weight_rom[71][38] = -32'd1944;
    weight_rom[71][39] = -32'd2255;
    weight_rom[71][40] = 32'd2632;
    weight_rom[71][41] = 32'd1046;
    weight_rom[71][42] = 32'd1575;
    weight_rom[71][43] = -32'd4871;
    weight_rom[71][44] = -32'd3246;
    weight_rom[71][45] = -32'd333;
    weight_rom[71][46] = 32'd4075;
    weight_rom[71][47] = -32'd3853;
    weight_rom[71][48] = 32'd3973;
    weight_rom[71][49] = 32'd4253;
    weight_rom[71][50] = 32'd4245;
    weight_rom[71][51] = 32'd1069;
    weight_rom[71][52] = -32'd5377;
    weight_rom[71][53] = -32'd2267;
    weight_rom[71][54] = 32'd4390;
    weight_rom[71][55] = 32'd5482;
    weight_rom[71][56] = -32'd864;
    weight_rom[71][57] = 32'd1037;
    weight_rom[71][58] = -32'd5526;
    weight_rom[71][59] = 32'd2498;
    weight_rom[71][60] = 32'd2465;
    weight_rom[71][61] = -32'd5966;
    weight_rom[71][62] = -32'd3180;
    weight_rom[71][63] = -32'd5720;
    weight_rom[72][0] = -32'd6481;
    weight_rom[72][1] = 32'd1861;
    weight_rom[72][2] = -32'd1053;
    weight_rom[72][3] = -32'd6404;
    weight_rom[72][4] = 32'd1748;
    weight_rom[72][5] = -32'd372;
    weight_rom[72][6] = -32'd6381;
    weight_rom[72][7] = 32'd870;
    weight_rom[72][8] = -32'd3663;
    weight_rom[72][9] = -32'd1052;
    weight_rom[72][10] = -32'd804;
    weight_rom[72][11] = 32'd4165;
    weight_rom[72][12] = -32'd3490;
    weight_rom[72][13] = -32'd658;
    weight_rom[72][14] = 32'd6352;
    weight_rom[72][15] = 32'd1444;
    weight_rom[72][16] = 32'd3979;
    weight_rom[72][17] = 32'd1297;
    weight_rom[72][18] = -32'd2538;
    weight_rom[72][19] = -32'd3925;
    weight_rom[72][20] = -32'd6496;
    weight_rom[72][21] = -32'd4622;
    weight_rom[72][22] = 32'd4074;
    weight_rom[72][23] = 32'd3050;
    weight_rom[72][24] = -32'd3029;
    weight_rom[72][25] = 32'd2928;
    weight_rom[72][26] = -32'd5672;
    weight_rom[72][27] = 32'd6131;
    weight_rom[72][28] = -32'd2091;
    weight_rom[72][29] = 32'd3945;
    weight_rom[72][30] = -32'd6469;
    weight_rom[72][31] = 32'd4798;
    weight_rom[72][32] = -32'd2425;
    weight_rom[72][33] = -32'd4673;
    weight_rom[72][34] = -32'd2420;
    weight_rom[72][35] = -32'd4537;
    weight_rom[72][36] = -32'd3007;
    weight_rom[72][37] = -32'd3316;
    weight_rom[72][38] = 32'd5368;
    weight_rom[72][39] = 32'd3108;
    weight_rom[72][40] = 32'd3477;
    weight_rom[72][41] = -32'd2850;
    weight_rom[72][42] = 32'd587;
    weight_rom[72][43] = 32'd1968;
    weight_rom[72][44] = 32'd5443;
    weight_rom[72][45] = 32'd4142;
    weight_rom[72][46] = -32'd1306;
    weight_rom[72][47] = 32'd2743;
    weight_rom[72][48] = -32'd4542;
    weight_rom[72][49] = -32'd1078;
    weight_rom[72][50] = 32'd1933;
    weight_rom[72][51] = 32'd438;
    weight_rom[72][52] = 32'd6049;
    weight_rom[72][53] = 32'd1677;
    weight_rom[72][54] = 32'd4489;
    weight_rom[72][55] = -32'd1205;
    weight_rom[72][56] = 32'd4186;
    weight_rom[72][57] = -32'd4075;
    weight_rom[72][58] = -32'd5602;
    weight_rom[72][59] = 32'd176;
    weight_rom[72][60] = -32'd4873;
    weight_rom[72][61] = -32'd5845;
    weight_rom[72][62] = 32'd2536;
    weight_rom[72][63] = -32'd1359;
    weight_rom[73][0] = 32'd4134;
    weight_rom[73][1] = -32'd5450;
    weight_rom[73][2] = -32'd3306;
    weight_rom[73][3] = -32'd410;
    weight_rom[73][4] = -32'd3405;
    weight_rom[73][5] = -32'd1155;
    weight_rom[73][6] = 32'd2143;
    weight_rom[73][7] = -32'd313;
    weight_rom[73][8] = -32'd4109;
    weight_rom[73][9] = 32'd1815;
    weight_rom[73][10] = 32'd2952;
    weight_rom[73][11] = -32'd4977;
    weight_rom[73][12] = 32'd524;
    weight_rom[73][13] = -32'd4002;
    weight_rom[73][14] = 32'd5732;
    weight_rom[73][15] = -32'd4779;
    weight_rom[73][16] = 32'd68;
    weight_rom[73][17] = -32'd5047;
    weight_rom[73][18] = 32'd3787;
    weight_rom[73][19] = -32'd5121;
    weight_rom[73][20] = -32'd4365;
    weight_rom[73][21] = -32'd6450;
    weight_rom[73][22] = 32'd4401;
    weight_rom[73][23] = -32'd1251;
    weight_rom[73][24] = -32'd1724;
    weight_rom[73][25] = 32'd467;
    weight_rom[73][26] = -32'd5309;
    weight_rom[73][27] = -32'd789;
    weight_rom[73][28] = 32'd138;
    weight_rom[73][29] = -32'd5184;
    weight_rom[73][30] = 32'd6269;
    weight_rom[73][31] = -32'd2759;
    weight_rom[73][32] = -32'd5286;
    weight_rom[73][33] = -32'd4568;
    weight_rom[73][34] = -32'd1400;
    weight_rom[73][35] = 32'd5061;
    weight_rom[73][36] = -32'd3292;
    weight_rom[73][37] = 32'd4713;
    weight_rom[73][38] = 32'd903;
    weight_rom[73][39] = -32'd6072;
    weight_rom[73][40] = 32'd5628;
    weight_rom[73][41] = -32'd2896;
    weight_rom[73][42] = -32'd4906;
    weight_rom[73][43] = 32'd6324;
    weight_rom[73][44] = -32'd3071;
    weight_rom[73][45] = -32'd890;
    weight_rom[73][46] = 32'd5860;
    weight_rom[73][47] = -32'd6276;
    weight_rom[73][48] = -32'd1749;
    weight_rom[73][49] = -32'd5595;
    weight_rom[73][50] = 32'd6146;
    weight_rom[73][51] = 32'd1263;
    weight_rom[73][52] = 32'd4027;
    weight_rom[73][53] = -32'd2946;
    weight_rom[73][54] = -32'd2579;
    weight_rom[73][55] = -32'd4046;
    weight_rom[73][56] = 32'd5316;
    weight_rom[73][57] = 32'd5254;
    weight_rom[73][58] = 32'd4591;
    weight_rom[73][59] = 32'd1974;
    weight_rom[73][60] = -32'd978;
    weight_rom[73][61] = -32'd560;
    weight_rom[73][62] = -32'd6033;
    weight_rom[73][63] = 32'd6079;
    weight_rom[74][0] = 32'd2711;
    weight_rom[74][1] = -32'd4435;
    weight_rom[74][2] = -32'd1887;
    weight_rom[74][3] = -32'd5815;
    weight_rom[74][4] = -32'd5559;
    weight_rom[74][5] = -32'd1980;
    weight_rom[74][6] = -32'd4220;
    weight_rom[74][7] = 32'd2145;
    weight_rom[74][8] = 32'd3664;
    weight_rom[74][9] = -32'd1342;
    weight_rom[74][10] = -32'd174;
    weight_rom[74][11] = 32'd583;
    weight_rom[74][12] = 32'd4981;
    weight_rom[74][13] = -32'd1733;
    weight_rom[74][14] = -32'd5987;
    weight_rom[74][15] = 32'd3294;
    weight_rom[74][16] = 32'd6122;
    weight_rom[74][17] = -32'd5323;
    weight_rom[74][18] = -32'd702;
    weight_rom[74][19] = 32'd4639;
    weight_rom[74][20] = 32'd2792;
    weight_rom[74][21] = 32'd1715;
    weight_rom[74][22] = -32'd2199;
    weight_rom[74][23] = -32'd5657;
    weight_rom[74][24] = 32'd5181;
    weight_rom[74][25] = 32'd4405;
    weight_rom[74][26] = 32'd6539;
    weight_rom[74][27] = -32'd2904;
    weight_rom[74][28] = 32'd1509;
    weight_rom[74][29] = 32'd1007;
    weight_rom[74][30] = 32'd6104;
    weight_rom[74][31] = -32'd423;
    weight_rom[74][32] = -32'd4235;
    weight_rom[74][33] = -32'd881;
    weight_rom[74][34] = -32'd3448;
    weight_rom[74][35] = -32'd543;
    weight_rom[74][36] = 32'd5794;
    weight_rom[74][37] = -32'd4340;
    weight_rom[74][38] = 32'd3436;
    weight_rom[74][39] = -32'd330;
    weight_rom[74][40] = -32'd3869;
    weight_rom[74][41] = -32'd1245;
    weight_rom[74][42] = -32'd2756;
    weight_rom[74][43] = 32'd5397;
    weight_rom[74][44] = 32'd5188;
    weight_rom[74][45] = 32'd3884;
    weight_rom[74][46] = -32'd1225;
    weight_rom[74][47] = -32'd1062;
    weight_rom[74][48] = -32'd1659;
    weight_rom[74][49] = -32'd2966;
    weight_rom[74][50] = 32'd2804;
    weight_rom[74][51] = -32'd1755;
    weight_rom[74][52] = -32'd529;
    weight_rom[74][53] = 32'd5368;
    weight_rom[74][54] = -32'd924;
    weight_rom[74][55] = 32'd224;
    weight_rom[74][56] = -32'd4983;
    weight_rom[74][57] = 32'd2283;
    weight_rom[74][58] = -32'd3763;
    weight_rom[74][59] = 32'd5107;
    weight_rom[74][60] = -32'd3313;
    weight_rom[74][61] = 32'd650;
    weight_rom[74][62] = 32'd4448;
    weight_rom[74][63] = 32'd510;
    weight_rom[75][0] = 32'd3001;
    weight_rom[75][1] = 32'd5223;
    weight_rom[75][2] = 32'd3379;
    weight_rom[75][3] = -32'd4996;
    weight_rom[75][4] = -32'd4864;
    weight_rom[75][5] = 32'd5629;
    weight_rom[75][6] = 32'd6043;
    weight_rom[75][7] = 32'd5725;
    weight_rom[75][8] = -32'd1964;
    weight_rom[75][9] = -32'd2959;
    weight_rom[75][10] = 32'd4894;
    weight_rom[75][11] = -32'd6478;
    weight_rom[75][12] = 32'd1977;
    weight_rom[75][13] = -32'd1125;
    weight_rom[75][14] = -32'd4393;
    weight_rom[75][15] = 32'd2057;
    weight_rom[75][16] = -32'd1077;
    weight_rom[75][17] = 32'd5369;
    weight_rom[75][18] = 32'd3910;
    weight_rom[75][19] = -32'd797;
    weight_rom[75][20] = 32'd2180;
    weight_rom[75][21] = -32'd685;
    weight_rom[75][22] = 32'd2537;
    weight_rom[75][23] = 32'd3719;
    weight_rom[75][24] = 32'd2181;
    weight_rom[75][25] = 32'd4212;
    weight_rom[75][26] = -32'd2272;
    weight_rom[75][27] = 32'd3909;
    weight_rom[75][28] = 32'd5381;
    weight_rom[75][29] = -32'd472;
    weight_rom[75][30] = -32'd1374;
    weight_rom[75][31] = 32'd1564;
    weight_rom[75][32] = 32'd6387;
    weight_rom[75][33] = 32'd1254;
    weight_rom[75][34] = -32'd5282;
    weight_rom[75][35] = 32'd846;
    weight_rom[75][36] = -32'd2644;
    weight_rom[75][37] = 32'd4639;
    weight_rom[75][38] = 32'd4086;
    weight_rom[75][39] = -32'd2145;
    weight_rom[75][40] = 32'd3905;
    weight_rom[75][41] = 32'd6537;
    weight_rom[75][42] = -32'd3424;
    weight_rom[75][43] = -32'd797;
    weight_rom[75][44] = -32'd5197;
    weight_rom[75][45] = 32'd1250;
    weight_rom[75][46] = 32'd3562;
    weight_rom[75][47] = 32'd3615;
    weight_rom[75][48] = -32'd4569;
    weight_rom[75][49] = 32'd6291;
    weight_rom[75][50] = 32'd5566;
    weight_rom[75][51] = 32'd4025;
    weight_rom[75][52] = -32'd3622;
    weight_rom[75][53] = 32'd1754;
    weight_rom[75][54] = -32'd383;
    weight_rom[75][55] = 32'd5348;
    weight_rom[75][56] = 32'd418;
    weight_rom[75][57] = 32'd1746;
    weight_rom[75][58] = 32'd2211;
    weight_rom[75][59] = -32'd780;
    weight_rom[75][60] = 32'd3255;
    weight_rom[75][61] = 32'd5083;
    weight_rom[75][62] = -32'd679;
    weight_rom[75][63] = -32'd2780;
    weight_rom[76][0] = 32'd3555;
    weight_rom[76][1] = 32'd1394;
    weight_rom[76][2] = -32'd6364;
    weight_rom[76][3] = -32'd5013;
    weight_rom[76][4] = -32'd4875;
    weight_rom[76][5] = 32'd4333;
    weight_rom[76][6] = -32'd4605;
    weight_rom[76][7] = 32'd3048;
    weight_rom[76][8] = -32'd5795;
    weight_rom[76][9] = 32'd6343;
    weight_rom[76][10] = 32'd5252;
    weight_rom[76][11] = -32'd2299;
    weight_rom[76][12] = 32'd432;
    weight_rom[76][13] = 32'd4293;
    weight_rom[76][14] = -32'd4826;
    weight_rom[76][15] = 32'd5984;
    weight_rom[76][16] = 32'd6345;
    weight_rom[76][17] = 32'd2217;
    weight_rom[76][18] = 32'd4226;
    weight_rom[76][19] = 32'd4547;
    weight_rom[76][20] = 32'd6108;
    weight_rom[76][21] = -32'd4793;
    weight_rom[76][22] = 32'd3553;
    weight_rom[76][23] = -32'd2808;
    weight_rom[76][24] = 32'd3766;
    weight_rom[76][25] = 32'd4500;
    weight_rom[76][26] = 32'd3253;
    weight_rom[76][27] = -32'd2277;
    weight_rom[76][28] = 32'd129;
    weight_rom[76][29] = -32'd4997;
    weight_rom[76][30] = 32'd2993;
    weight_rom[76][31] = -32'd1164;
    weight_rom[76][32] = -32'd732;
    weight_rom[76][33] = -32'd5496;
    weight_rom[76][34] = -32'd4207;
    weight_rom[76][35] = 32'd2136;
    weight_rom[76][36] = 32'd3611;
    weight_rom[76][37] = -32'd6380;
    weight_rom[76][38] = -32'd2072;
    weight_rom[76][39] = 32'd5512;
    weight_rom[76][40] = 32'd3126;
    weight_rom[76][41] = -32'd5833;
    weight_rom[76][42] = -32'd3754;
    weight_rom[76][43] = -32'd6029;
    weight_rom[76][44] = 32'd2052;
    weight_rom[76][45] = 32'd5067;
    weight_rom[76][46] = -32'd211;
    weight_rom[76][47] = -32'd2113;
    weight_rom[76][48] = 32'd3911;
    weight_rom[76][49] = 32'd1261;
    weight_rom[76][50] = 32'd224;
    weight_rom[76][51] = 32'd305;
    weight_rom[76][52] = 32'd5681;
    weight_rom[76][53] = -32'd5611;
    weight_rom[76][54] = -32'd4490;
    weight_rom[76][55] = 32'd3989;
    weight_rom[76][56] = -32'd2824;
    weight_rom[76][57] = -32'd5249;
    weight_rom[76][58] = 32'd562;
    weight_rom[76][59] = 32'd5258;
    weight_rom[76][60] = -32'd3119;
    weight_rom[76][61] = -32'd5181;
    weight_rom[76][62] = 32'd1791;
    weight_rom[76][63] = -32'd4977;
    weight_rom[77][0] = -32'd5583;
    weight_rom[77][1] = -32'd6433;
    weight_rom[77][2] = -32'd5032;
    weight_rom[77][3] = 32'd1955;
    weight_rom[77][4] = -32'd4562;
    weight_rom[77][5] = 32'd6095;
    weight_rom[77][6] = -32'd1119;
    weight_rom[77][7] = -32'd3736;
    weight_rom[77][8] = 32'd6148;
    weight_rom[77][9] = -32'd1188;
    weight_rom[77][10] = -32'd1026;
    weight_rom[77][11] = -32'd1750;
    weight_rom[77][12] = -32'd2302;
    weight_rom[77][13] = 32'd3062;
    weight_rom[77][14] = 32'd2961;
    weight_rom[77][15] = -32'd5649;
    weight_rom[77][16] = 32'd2200;
    weight_rom[77][17] = 32'd4316;
    weight_rom[77][18] = 32'd4686;
    weight_rom[77][19] = 32'd5152;
    weight_rom[77][20] = 32'd3421;
    weight_rom[77][21] = 32'd6002;
    weight_rom[77][22] = 32'd2027;
    weight_rom[77][23] = -32'd881;
    weight_rom[77][24] = -32'd598;
    weight_rom[77][25] = -32'd195;
    weight_rom[77][26] = 32'd4019;
    weight_rom[77][27] = -32'd2629;
    weight_rom[77][28] = 32'd16;
    weight_rom[77][29] = 32'd6298;
    weight_rom[77][30] = -32'd2021;
    weight_rom[77][31] = -32'd950;
    weight_rom[77][32] = 32'd417;
    weight_rom[77][33] = 32'd5761;
    weight_rom[77][34] = 32'd3899;
    weight_rom[77][35] = 32'd2347;
    weight_rom[77][36] = -32'd1400;
    weight_rom[77][37] = 32'd154;
    weight_rom[77][38] = -32'd869;
    weight_rom[77][39] = -32'd6396;
    weight_rom[77][40] = -32'd5717;
    weight_rom[77][41] = 32'd1029;
    weight_rom[77][42] = -32'd1164;
    weight_rom[77][43] = -32'd1804;
    weight_rom[77][44] = 32'd5334;
    weight_rom[77][45] = -32'd1167;
    weight_rom[77][46] = 32'd5210;
    weight_rom[77][47] = 32'd835;
    weight_rom[77][48] = 32'd2716;
    weight_rom[77][49] = 32'd2749;
    weight_rom[77][50] = -32'd5019;
    weight_rom[77][51] = -32'd5023;
    weight_rom[77][52] = -32'd2036;
    weight_rom[77][53] = 32'd5360;
    weight_rom[77][54] = -32'd6146;
    weight_rom[77][55] = -32'd5690;
    weight_rom[77][56] = -32'd5936;
    weight_rom[77][57] = 32'd1365;
    weight_rom[77][58] = 32'd4363;
    weight_rom[77][59] = 32'd3285;
    weight_rom[77][60] = 32'd5003;
    weight_rom[77][61] = 32'd4229;
    weight_rom[77][62] = -32'd3653;
    weight_rom[77][63] = 32'd2667;
    weight_rom[78][0] = -32'd1855;
    weight_rom[78][1] = -32'd5223;
    weight_rom[78][2] = -32'd5950;
    weight_rom[78][3] = 32'd3224;
    weight_rom[78][4] = -32'd4733;
    weight_rom[78][5] = -32'd4924;
    weight_rom[78][6] = -32'd5434;
    weight_rom[78][7] = -32'd6144;
    weight_rom[78][8] = 32'd5030;
    weight_rom[78][9] = 32'd5165;
    weight_rom[78][10] = -32'd2925;
    weight_rom[78][11] = -32'd1360;
    weight_rom[78][12] = -32'd2188;
    weight_rom[78][13] = 32'd3529;
    weight_rom[78][14] = 32'd4165;
    weight_rom[78][15] = -32'd5805;
    weight_rom[78][16] = 32'd1765;
    weight_rom[78][17] = 32'd4967;
    weight_rom[78][18] = 32'd5460;
    weight_rom[78][19] = -32'd5734;
    weight_rom[78][20] = 32'd5908;
    weight_rom[78][21] = 32'd388;
    weight_rom[78][22] = -32'd4566;
    weight_rom[78][23] = 32'd2430;
    weight_rom[78][24] = 32'd1707;
    weight_rom[78][25] = -32'd2180;
    weight_rom[78][26] = 32'd4692;
    weight_rom[78][27] = -32'd3506;
    weight_rom[78][28] = -32'd5895;
    weight_rom[78][29] = -32'd3739;
    weight_rom[78][30] = 32'd2242;
    weight_rom[78][31] = -32'd2224;
    weight_rom[78][32] = 32'd4897;
    weight_rom[78][33] = 32'd3344;
    weight_rom[78][34] = 32'd2327;
    weight_rom[78][35] = 32'd5658;
    weight_rom[78][36] = -32'd4728;
    weight_rom[78][37] = 32'd3531;
    weight_rom[78][38] = 32'd4567;
    weight_rom[78][39] = 32'd692;
    weight_rom[78][40] = -32'd1478;
    weight_rom[78][41] = -32'd5471;
    weight_rom[78][42] = 32'd2674;
    weight_rom[78][43] = 32'd4278;
    weight_rom[78][44] = -32'd4341;
    weight_rom[78][45] = 32'd1367;
    weight_rom[78][46] = 32'd5344;
    weight_rom[78][47] = -32'd3866;
    weight_rom[78][48] = -32'd4058;
    weight_rom[78][49] = -32'd6457;
    weight_rom[78][50] = 32'd369;
    weight_rom[78][51] = -32'd4861;
    weight_rom[78][52] = -32'd4443;
    weight_rom[78][53] = 32'd6000;
    weight_rom[78][54] = 32'd5857;
    weight_rom[78][55] = 32'd2524;
    weight_rom[78][56] = 32'd2209;
    weight_rom[78][57] = -32'd4968;
    weight_rom[78][58] = -32'd4914;
    weight_rom[78][59] = -32'd149;
    weight_rom[78][60] = 32'd5135;
    weight_rom[78][61] = -32'd3800;
    weight_rom[78][62] = 32'd2320;
    weight_rom[78][63] = 32'd1898;
    weight_rom[79][0] = -32'd5034;
    weight_rom[79][1] = 32'd2143;
    weight_rom[79][2] = -32'd6019;
    weight_rom[79][3] = 32'd1092;
    weight_rom[79][4] = 32'd1846;
    weight_rom[79][5] = 32'd3025;
    weight_rom[79][6] = 32'd6512;
    weight_rom[79][7] = -32'd3116;
    weight_rom[79][8] = 32'd5606;
    weight_rom[79][9] = -32'd3539;
    weight_rom[79][10] = 32'd1210;
    weight_rom[79][11] = 32'd2561;
    weight_rom[79][12] = 32'd2221;
    weight_rom[79][13] = -32'd6409;
    weight_rom[79][14] = -32'd3755;
    weight_rom[79][15] = -32'd2854;
    weight_rom[79][16] = -32'd4378;
    weight_rom[79][17] = 32'd940;
    weight_rom[79][18] = -32'd904;
    weight_rom[79][19] = 32'd5026;
    weight_rom[79][20] = 32'd2654;
    weight_rom[79][21] = -32'd3383;
    weight_rom[79][22] = 32'd4926;
    weight_rom[79][23] = -32'd2196;
    weight_rom[79][24] = -32'd3297;
    weight_rom[79][25] = 32'd3821;
    weight_rom[79][26] = 32'd6522;
    weight_rom[79][27] = -32'd4853;
    weight_rom[79][28] = -32'd6096;
    weight_rom[79][29] = -32'd5672;
    weight_rom[79][30] = 32'd4003;
    weight_rom[79][31] = 32'd841;
    weight_rom[79][32] = 32'd6495;
    weight_rom[79][33] = 32'd1135;
    weight_rom[79][34] = 32'd615;
    weight_rom[79][35] = 32'd6513;
    weight_rom[79][36] = -32'd6413;
    weight_rom[79][37] = 32'd5698;
    weight_rom[79][38] = -32'd1792;
    weight_rom[79][39] = 32'd3154;
    weight_rom[79][40] = -32'd2847;
    weight_rom[79][41] = -32'd4528;
    weight_rom[79][42] = -32'd3703;
    weight_rom[79][43] = 32'd2641;
    weight_rom[79][44] = 32'd6138;
    weight_rom[79][45] = 32'd1704;
    weight_rom[79][46] = -32'd5407;
    weight_rom[79][47] = 32'd3171;
    weight_rom[79][48] = -32'd1746;
    weight_rom[79][49] = 32'd238;
    weight_rom[79][50] = -32'd4890;
    weight_rom[79][51] = 32'd483;
    weight_rom[79][52] = 32'd827;
    weight_rom[79][53] = -32'd5535;
    weight_rom[79][54] = -32'd3398;
    weight_rom[79][55] = 32'd942;
    weight_rom[79][56] = 32'd4754;
    weight_rom[79][57] = -32'd5522;
    weight_rom[79][58] = -32'd4852;
    weight_rom[79][59] = 32'd1352;
    weight_rom[79][60] = -32'd3978;
    weight_rom[79][61] = -32'd1388;
    weight_rom[79][62] = 32'd3568;
    weight_rom[79][63] = -32'd1652;
    weight_rom[80][0] = 32'd4759;
    weight_rom[80][1] = -32'd6487;
    weight_rom[80][2] = 32'd4659;
    weight_rom[80][3] = 32'd6057;
    weight_rom[80][4] = -32'd4169;
    weight_rom[80][5] = 32'd5745;
    weight_rom[80][6] = 32'd28;
    weight_rom[80][7] = 32'd1246;
    weight_rom[80][8] = 32'd6486;
    weight_rom[80][9] = -32'd3760;
    weight_rom[80][10] = 32'd5404;
    weight_rom[80][11] = -32'd1460;
    weight_rom[80][12] = 32'd6476;
    weight_rom[80][13] = -32'd1098;
    weight_rom[80][14] = 32'd76;
    weight_rom[80][15] = -32'd3123;
    weight_rom[80][16] = 32'd5006;
    weight_rom[80][17] = 32'd228;
    weight_rom[80][18] = -32'd2374;
    weight_rom[80][19] = -32'd677;
    weight_rom[80][20] = -32'd2646;
    weight_rom[80][21] = 32'd7;
    weight_rom[80][22] = 32'd512;
    weight_rom[80][23] = -32'd5811;
    weight_rom[80][24] = 32'd2693;
    weight_rom[80][25] = -32'd638;
    weight_rom[80][26] = -32'd3388;
    weight_rom[80][27] = -32'd3192;
    weight_rom[80][28] = 32'd670;
    weight_rom[80][29] = 32'd1243;
    weight_rom[80][30] = 32'd5855;
    weight_rom[80][31] = 32'd4595;
    weight_rom[80][32] = 32'd1084;
    weight_rom[80][33] = 32'd4304;
    weight_rom[80][34] = -32'd326;
    weight_rom[80][35] = 32'd2885;
    weight_rom[80][36] = 32'd580;
    weight_rom[80][37] = 32'd5363;
    weight_rom[80][38] = 32'd3852;
    weight_rom[80][39] = -32'd196;
    weight_rom[80][40] = -32'd2562;
    weight_rom[80][41] = -32'd792;
    weight_rom[80][42] = -32'd1747;
    weight_rom[80][43] = -32'd532;
    weight_rom[80][44] = -32'd617;
    weight_rom[80][45] = -32'd1082;
    weight_rom[80][46] = 32'd5721;
    weight_rom[80][47] = -32'd5868;
    weight_rom[80][48] = -32'd5166;
    weight_rom[80][49] = -32'd6061;
    weight_rom[80][50] = 32'd1212;
    weight_rom[80][51] = 32'd5722;
    weight_rom[80][52] = 32'd5816;
    weight_rom[80][53] = 32'd424;
    weight_rom[80][54] = -32'd3408;
    weight_rom[80][55] = 32'd5340;
    weight_rom[80][56] = -32'd4418;
    weight_rom[80][57] = 32'd357;
    weight_rom[80][58] = 32'd744;
    weight_rom[80][59] = -32'd2286;
    weight_rom[80][60] = 32'd1492;
    weight_rom[80][61] = -32'd2403;
    weight_rom[80][62] = -32'd351;
    weight_rom[80][63] = 32'd5910;
    weight_rom[81][0] = 32'd1616;
    weight_rom[81][1] = -32'd4445;
    weight_rom[81][2] = 32'd2669;
    weight_rom[81][3] = -32'd1640;
    weight_rom[81][4] = -32'd2022;
    weight_rom[81][5] = -32'd4178;
    weight_rom[81][6] = 32'd1250;
    weight_rom[81][7] = -32'd5879;
    weight_rom[81][8] = -32'd4274;
    weight_rom[81][9] = -32'd6145;
    weight_rom[81][10] = -32'd3792;
    weight_rom[81][11] = -32'd672;
    weight_rom[81][12] = 32'd2121;
    weight_rom[81][13] = -32'd244;
    weight_rom[81][14] = 32'd4465;
    weight_rom[81][15] = -32'd3316;
    weight_rom[81][16] = -32'd950;
    weight_rom[81][17] = -32'd911;
    weight_rom[81][18] = 32'd1077;
    weight_rom[81][19] = 32'd136;
    weight_rom[81][20] = -32'd5172;
    weight_rom[81][21] = 32'd2354;
    weight_rom[81][22] = -32'd2851;
    weight_rom[81][23] = -32'd1652;
    weight_rom[81][24] = -32'd948;
    weight_rom[81][25] = -32'd4149;
    weight_rom[81][26] = -32'd6024;
    weight_rom[81][27] = -32'd1896;
    weight_rom[81][28] = -32'd810;
    weight_rom[81][29] = 32'd3130;
    weight_rom[81][30] = -32'd1307;
    weight_rom[81][31] = -32'd3912;
    weight_rom[81][32] = 32'd4095;
    weight_rom[81][33] = -32'd5502;
    weight_rom[81][34] = 32'd5536;
    weight_rom[81][35] = -32'd2788;
    weight_rom[81][36] = 32'd6236;
    weight_rom[81][37] = 32'd4189;
    weight_rom[81][38] = 32'd5780;
    weight_rom[81][39] = -32'd5434;
    weight_rom[81][40] = 32'd6330;
    weight_rom[81][41] = 32'd137;
    weight_rom[81][42] = -32'd1429;
    weight_rom[81][43] = -32'd5831;
    weight_rom[81][44] = 32'd5842;
    weight_rom[81][45] = -32'd4662;
    weight_rom[81][46] = 32'd4266;
    weight_rom[81][47] = 32'd4620;
    weight_rom[81][48] = 32'd1680;
    weight_rom[81][49] = 32'd907;
    weight_rom[81][50] = -32'd229;
    weight_rom[81][51] = -32'd2511;
    weight_rom[81][52] = -32'd6503;
    weight_rom[81][53] = -32'd2577;
    weight_rom[81][54] = -32'd5460;
    weight_rom[81][55] = -32'd4948;
    weight_rom[81][56] = 32'd4094;
    weight_rom[81][57] = -32'd1274;
    weight_rom[81][58] = 32'd5850;
    weight_rom[81][59] = 32'd6338;
    weight_rom[81][60] = -32'd5403;
    weight_rom[81][61] = -32'd1308;
    weight_rom[81][62] = 32'd1543;
    weight_rom[81][63] = -32'd6262;
    weight_rom[82][0] = -32'd2216;
    weight_rom[82][1] = 32'd638;
    weight_rom[82][2] = -32'd338;
    weight_rom[82][3] = -32'd2808;
    weight_rom[82][4] = 32'd5200;
    weight_rom[82][5] = -32'd5682;
    weight_rom[82][6] = -32'd5674;
    weight_rom[82][7] = -32'd47;
    weight_rom[82][8] = -32'd1360;
    weight_rom[82][9] = 32'd1987;
    weight_rom[82][10] = 32'd1611;
    weight_rom[82][11] = -32'd3440;
    weight_rom[82][12] = 32'd757;
    weight_rom[82][13] = -32'd6302;
    weight_rom[82][14] = 32'd3051;
    weight_rom[82][15] = 32'd5324;
    weight_rom[82][16] = -32'd4427;
    weight_rom[82][17] = -32'd2399;
    weight_rom[82][18] = -32'd1688;
    weight_rom[82][19] = 32'd1659;
    weight_rom[82][20] = 32'd3693;
    weight_rom[82][21] = -32'd5554;
    weight_rom[82][22] = -32'd980;
    weight_rom[82][23] = 32'd5825;
    weight_rom[82][24] = -32'd753;
    weight_rom[82][25] = 32'd4652;
    weight_rom[82][26] = -32'd1164;
    weight_rom[82][27] = 32'd2280;
    weight_rom[82][28] = 32'd4445;
    weight_rom[82][29] = -32'd6128;
    weight_rom[82][30] = 32'd3713;
    weight_rom[82][31] = 32'd5694;
    weight_rom[82][32] = -32'd2268;
    weight_rom[82][33] = -32'd303;
    weight_rom[82][34] = -32'd5600;
    weight_rom[82][35] = 32'd4977;
    weight_rom[82][36] = -32'd1715;
    weight_rom[82][37] = 32'd5088;
    weight_rom[82][38] = 32'd1614;
    weight_rom[82][39] = 32'd6192;
    weight_rom[82][40] = 32'd1871;
    weight_rom[82][41] = -32'd3161;
    weight_rom[82][42] = 32'd6244;
    weight_rom[82][43] = -32'd958;
    weight_rom[82][44] = 32'd2317;
    weight_rom[82][45] = -32'd5327;
    weight_rom[82][46] = 32'd3818;
    weight_rom[82][47] = -32'd3955;
    weight_rom[82][48] = -32'd4962;
    weight_rom[82][49] = 32'd5515;
    weight_rom[82][50] = 32'd1606;
    weight_rom[82][51] = 32'd4843;
    weight_rom[82][52] = -32'd3432;
    weight_rom[82][53] = -32'd1404;
    weight_rom[82][54] = 32'd5616;
    weight_rom[82][55] = 32'd446;
    weight_rom[82][56] = 32'd4632;
    weight_rom[82][57] = 32'd1164;
    weight_rom[82][58] = -32'd1114;
    weight_rom[82][59] = 32'd2193;
    weight_rom[82][60] = -32'd1421;
    weight_rom[82][61] = -32'd4581;
    weight_rom[82][62] = -32'd572;
    weight_rom[82][63] = -32'd2572;
    weight_rom[83][0] = -32'd5720;
    weight_rom[83][1] = 32'd2515;
    weight_rom[83][2] = -32'd5271;
    weight_rom[83][3] = 32'd4831;
    weight_rom[83][4] = -32'd341;
    weight_rom[83][5] = 32'd3160;
    weight_rom[83][6] = 32'd3276;
    weight_rom[83][7] = 32'd1269;
    weight_rom[83][8] = 32'd3384;
    weight_rom[83][9] = -32'd1723;
    weight_rom[83][10] = 32'd1724;
    weight_rom[83][11] = -32'd1661;
    weight_rom[83][12] = 32'd3023;
    weight_rom[83][13] = -32'd3148;
    weight_rom[83][14] = 32'd553;
    weight_rom[83][15] = -32'd3282;
    weight_rom[83][16] = -32'd6388;
    weight_rom[83][17] = -32'd857;
    weight_rom[83][18] = 32'd1324;
    weight_rom[83][19] = 32'd5588;
    weight_rom[83][20] = 32'd1889;
    weight_rom[83][21] = -32'd2952;
    weight_rom[83][22] = -32'd6061;
    weight_rom[83][23] = 32'd1857;
    weight_rom[83][24] = 32'd1957;
    weight_rom[83][25] = 32'd5014;
    weight_rom[83][26] = -32'd4848;
    weight_rom[83][27] = -32'd5733;
    weight_rom[83][28] = -32'd4447;
    weight_rom[83][29] = 32'd2080;
    weight_rom[83][30] = -32'd3068;
    weight_rom[83][31] = 32'd2478;
    weight_rom[83][32] = -32'd2546;
    weight_rom[83][33] = 32'd1705;
    weight_rom[83][34] = -32'd2875;
    weight_rom[83][35] = -32'd5908;
    weight_rom[83][36] = -32'd1871;
    weight_rom[83][37] = -32'd3942;
    weight_rom[83][38] = 32'd3167;
    weight_rom[83][39] = 32'd236;
    weight_rom[83][40] = 32'd2853;
    weight_rom[83][41] = -32'd2405;
    weight_rom[83][42] = 32'd5959;
    weight_rom[83][43] = -32'd405;
    weight_rom[83][44] = -32'd2600;
    weight_rom[83][45] = -32'd6335;
    weight_rom[83][46] = -32'd3920;
    weight_rom[83][47] = 32'd4907;
    weight_rom[83][48] = 32'd6369;
    weight_rom[83][49] = 32'd6139;
    weight_rom[83][50] = -32'd6421;
    weight_rom[83][51] = 32'd3461;
    weight_rom[83][52] = 32'd5746;
    weight_rom[83][53] = -32'd4198;
    weight_rom[83][54] = 32'd1045;
    weight_rom[83][55] = 32'd4973;
    weight_rom[83][56] = 32'd5430;
    weight_rom[83][57] = -32'd5384;
    weight_rom[83][58] = -32'd2268;
    weight_rom[83][59] = -32'd5978;
    weight_rom[83][60] = 32'd2796;
    weight_rom[83][61] = 32'd46;
    weight_rom[83][62] = 32'd5165;
    weight_rom[83][63] = 32'd5519;
    weight_rom[84][0] = -32'd2477;
    weight_rom[84][1] = 32'd1991;
    weight_rom[84][2] = -32'd109;
    weight_rom[84][3] = -32'd3622;
    weight_rom[84][4] = 32'd2196;
    weight_rom[84][5] = 32'd976;
    weight_rom[84][6] = -32'd3802;
    weight_rom[84][7] = -32'd2172;
    weight_rom[84][8] = 32'd2569;
    weight_rom[84][9] = 32'd4775;
    weight_rom[84][10] = 32'd3055;
    weight_rom[84][11] = -32'd3574;
    weight_rom[84][12] = -32'd456;
    weight_rom[84][13] = 32'd3411;
    weight_rom[84][14] = 32'd1184;
    weight_rom[84][15] = -32'd2989;
    weight_rom[84][16] = 32'd783;
    weight_rom[84][17] = 32'd3589;
    weight_rom[84][18] = 32'd2694;
    weight_rom[84][19] = -32'd6303;
    weight_rom[84][20] = -32'd5922;
    weight_rom[84][21] = 32'd4023;
    weight_rom[84][22] = -32'd4877;
    weight_rom[84][23] = 32'd2247;
    weight_rom[84][24] = 32'd5718;
    weight_rom[84][25] = -32'd441;
    weight_rom[84][26] = -32'd6259;
    weight_rom[84][27] = -32'd3794;
    weight_rom[84][28] = -32'd6226;
    weight_rom[84][29] = 32'd423;
    weight_rom[84][30] = 32'd6426;
    weight_rom[84][31] = 32'd4237;
    weight_rom[84][32] = -32'd1275;
    weight_rom[84][33] = 32'd4307;
    weight_rom[84][34] = -32'd1966;
    weight_rom[84][35] = -32'd3524;
    weight_rom[84][36] = -32'd2043;
    weight_rom[84][37] = -32'd2828;
    weight_rom[84][38] = 32'd3998;
    weight_rom[84][39] = 32'd1496;
    weight_rom[84][40] = 32'd6247;
    weight_rom[84][41] = -32'd5413;
    weight_rom[84][42] = 32'd3933;
    weight_rom[84][43] = 32'd5617;
    weight_rom[84][44] = -32'd4085;
    weight_rom[84][45] = 32'd4895;
    weight_rom[84][46] = 32'd3999;
    weight_rom[84][47] = -32'd1932;
    weight_rom[84][48] = 32'd3678;
    weight_rom[84][49] = 32'd531;
    weight_rom[84][50] = -32'd3999;
    weight_rom[84][51] = -32'd3305;
    weight_rom[84][52] = -32'd4311;
    weight_rom[84][53] = 32'd1023;
    weight_rom[84][54] = 32'd2189;
    weight_rom[84][55] = -32'd1179;
    weight_rom[84][56] = -32'd3076;
    weight_rom[84][57] = -32'd904;
    weight_rom[84][58] = 32'd1398;
    weight_rom[84][59] = -32'd2272;
    weight_rom[84][60] = 32'd2089;
    weight_rom[84][61] = 32'd3953;
    weight_rom[84][62] = -32'd27;
    weight_rom[84][63] = -32'd2347;
    weight_rom[85][0] = -32'd2291;
    weight_rom[85][1] = -32'd3614;
    weight_rom[85][2] = -32'd347;
    weight_rom[85][3] = 32'd6071;
    weight_rom[85][4] = -32'd4294;
    weight_rom[85][5] = 32'd4480;
    weight_rom[85][6] = 32'd5217;
    weight_rom[85][7] = 32'd3550;
    weight_rom[85][8] = -32'd4536;
    weight_rom[85][9] = -32'd351;
    weight_rom[85][10] = -32'd4829;
    weight_rom[85][11] = -32'd5594;
    weight_rom[85][12] = -32'd5765;
    weight_rom[85][13] = -32'd4756;
    weight_rom[85][14] = 32'd109;
    weight_rom[85][15] = 32'd3400;
    weight_rom[85][16] = 32'd359;
    weight_rom[85][17] = 32'd1335;
    weight_rom[85][18] = 32'd2469;
    weight_rom[85][19] = -32'd303;
    weight_rom[85][20] = -32'd1834;
    weight_rom[85][21] = -32'd528;
    weight_rom[85][22] = 32'd3480;
    weight_rom[85][23] = 32'd1733;
    weight_rom[85][24] = -32'd5714;
    weight_rom[85][25] = -32'd5561;
    weight_rom[85][26] = -32'd1829;
    weight_rom[85][27] = 32'd4050;
    weight_rom[85][28] = -32'd667;
    weight_rom[85][29] = -32'd5200;
    weight_rom[85][30] = -32'd6215;
    weight_rom[85][31] = 32'd736;
    weight_rom[85][32] = 32'd2261;
    weight_rom[85][33] = 32'd3715;
    weight_rom[85][34] = 32'd3701;
    weight_rom[85][35] = 32'd5208;
    weight_rom[85][36] = 32'd269;
    weight_rom[85][37] = -32'd2766;
    weight_rom[85][38] = 32'd4522;
    weight_rom[85][39] = -32'd3452;
    weight_rom[85][40] = -32'd1609;
    weight_rom[85][41] = -32'd2579;
    weight_rom[85][42] = -32'd3386;
    weight_rom[85][43] = 32'd1849;
    weight_rom[85][44] = -32'd2572;
    weight_rom[85][45] = -32'd3454;
    weight_rom[85][46] = 32'd4589;
    weight_rom[85][47] = 32'd2918;
    weight_rom[85][48] = -32'd1438;
    weight_rom[85][49] = -32'd547;
    weight_rom[85][50] = -32'd113;
    weight_rom[85][51] = -32'd6077;
    weight_rom[85][52] = -32'd5069;
    weight_rom[85][53] = 32'd6002;
    weight_rom[85][54] = 32'd5394;
    weight_rom[85][55] = -32'd235;
    weight_rom[85][56] = 32'd5294;
    weight_rom[85][57] = -32'd4262;
    weight_rom[85][58] = 32'd5641;
    weight_rom[85][59] = 32'd1616;
    weight_rom[85][60] = 32'd1634;
    weight_rom[85][61] = -32'd766;
    weight_rom[85][62] = 32'd4480;
    weight_rom[85][63] = -32'd3247;
    weight_rom[86][0] = 32'd3009;
    weight_rom[86][1] = 32'd2781;
    weight_rom[86][2] = -32'd4283;
    weight_rom[86][3] = -32'd6394;
    weight_rom[86][4] = -32'd4033;
    weight_rom[86][5] = -32'd4721;
    weight_rom[86][6] = -32'd3864;
    weight_rom[86][7] = -32'd5156;
    weight_rom[86][8] = 32'd4139;
    weight_rom[86][9] = 32'd6136;
    weight_rom[86][10] = 32'd2828;
    weight_rom[86][11] = 32'd1355;
    weight_rom[86][12] = 32'd816;
    weight_rom[86][13] = 32'd462;
    weight_rom[86][14] = -32'd2653;
    weight_rom[86][15] = -32'd658;
    weight_rom[86][16] = 32'd2875;
    weight_rom[86][17] = 32'd5144;
    weight_rom[86][18] = -32'd1644;
    weight_rom[86][19] = 32'd2460;
    weight_rom[86][20] = 32'd5987;
    weight_rom[86][21] = 32'd610;
    weight_rom[86][22] = -32'd6553;
    weight_rom[86][23] = -32'd3945;
    weight_rom[86][24] = 32'd4256;
    weight_rom[86][25] = -32'd1470;
    weight_rom[86][26] = 32'd3719;
    weight_rom[86][27] = -32'd4627;
    weight_rom[86][28] = -32'd3440;
    weight_rom[86][29] = -32'd4292;
    weight_rom[86][30] = 32'd1356;
    weight_rom[86][31] = 32'd3663;
    weight_rom[86][32] = 32'd2388;
    weight_rom[86][33] = -32'd2921;
    weight_rom[86][34] = 32'd6455;
    weight_rom[86][35] = -32'd3195;
    weight_rom[86][36] = -32'd777;
    weight_rom[86][37] = -32'd1611;
    weight_rom[86][38] = -32'd1375;
    weight_rom[86][39] = -32'd216;
    weight_rom[86][40] = 32'd3956;
    weight_rom[86][41] = 32'd6115;
    weight_rom[86][42] = -32'd5661;
    weight_rom[86][43] = -32'd2468;
    weight_rom[86][44] = -32'd5334;
    weight_rom[86][45] = -32'd3781;
    weight_rom[86][46] = -32'd2763;
    weight_rom[86][47] = -32'd2369;
    weight_rom[86][48] = 32'd1029;
    weight_rom[86][49] = 32'd5832;
    weight_rom[86][50] = 32'd5904;
    weight_rom[86][51] = -32'd5218;
    weight_rom[86][52] = 32'd919;
    weight_rom[86][53] = 32'd40;
    weight_rom[86][54] = -32'd2023;
    weight_rom[86][55] = -32'd5630;
    weight_rom[86][56] = -32'd2350;
    weight_rom[86][57] = 32'd6384;
    weight_rom[86][58] = 32'd4416;
    weight_rom[86][59] = -32'd5815;
    weight_rom[86][60] = -32'd2850;
    weight_rom[86][61] = -32'd123;
    weight_rom[86][62] = 32'd3949;
    weight_rom[86][63] = 32'd448;
    weight_rom[87][0] = 32'd1802;
    weight_rom[87][1] = -32'd3443;
    weight_rom[87][2] = -32'd867;
    weight_rom[87][3] = 32'd6158;
    weight_rom[87][4] = -32'd6017;
    weight_rom[87][5] = 32'd3870;
    weight_rom[87][6] = -32'd4054;
    weight_rom[87][7] = -32'd5568;
    weight_rom[87][8] = -32'd3611;
    weight_rom[87][9] = -32'd4121;
    weight_rom[87][10] = 32'd5361;
    weight_rom[87][11] = 32'd2204;
    weight_rom[87][12] = 32'd5998;
    weight_rom[87][13] = -32'd3732;
    weight_rom[87][14] = 32'd852;
    weight_rom[87][15] = 32'd3626;
    weight_rom[87][16] = 32'd5115;
    weight_rom[87][17] = -32'd742;
    weight_rom[87][18] = -32'd4366;
    weight_rom[87][19] = 32'd2919;
    weight_rom[87][20] = 32'd5;
    weight_rom[87][21] = -32'd880;
    weight_rom[87][22] = -32'd1093;
    weight_rom[87][23] = -32'd1070;
    weight_rom[87][24] = -32'd2721;
    weight_rom[87][25] = 32'd3978;
    weight_rom[87][26] = 32'd867;
    weight_rom[87][27] = -32'd2062;
    weight_rom[87][28] = -32'd5903;
    weight_rom[87][29] = 32'd890;
    weight_rom[87][30] = 32'd2090;
    weight_rom[87][31] = -32'd6341;
    weight_rom[87][32] = -32'd2421;
    weight_rom[87][33] = 32'd5778;
    weight_rom[87][34] = -32'd3399;
    weight_rom[87][35] = -32'd3661;
    weight_rom[87][36] = 32'd4979;
    weight_rom[87][37] = -32'd1398;
    weight_rom[87][38] = -32'd5881;
    weight_rom[87][39] = -32'd928;
    weight_rom[87][40] = -32'd858;
    weight_rom[87][41] = 32'd5828;
    weight_rom[87][42] = -32'd2399;
    weight_rom[87][43] = 32'd331;
    weight_rom[87][44] = -32'd4667;
    weight_rom[87][45] = 32'd3093;
    weight_rom[87][46] = 32'd5927;
    weight_rom[87][47] = 32'd5320;
    weight_rom[87][48] = 32'd5391;
    weight_rom[87][49] = 32'd2275;
    weight_rom[87][50] = -32'd1525;
    weight_rom[87][51] = 32'd2994;
    weight_rom[87][52] = 32'd4742;
    weight_rom[87][53] = -32'd5466;
    weight_rom[87][54] = 32'd1592;
    weight_rom[87][55] = -32'd2907;
    weight_rom[87][56] = 32'd686;
    weight_rom[87][57] = 32'd801;
    weight_rom[87][58] = 32'd6494;
    weight_rom[87][59] = -32'd6240;
    weight_rom[87][60] = -32'd1598;
    weight_rom[87][61] = 32'd4571;
    weight_rom[87][62] = -32'd1173;
    weight_rom[87][63] = 32'd4244;
    weight_rom[88][0] = 32'd5075;
    weight_rom[88][1] = -32'd2288;
    weight_rom[88][2] = -32'd1330;
    weight_rom[88][3] = -32'd5987;
    weight_rom[88][4] = -32'd4339;
    weight_rom[88][5] = -32'd3910;
    weight_rom[88][6] = -32'd6074;
    weight_rom[88][7] = 32'd2990;
    weight_rom[88][8] = -32'd3619;
    weight_rom[88][9] = 32'd4831;
    weight_rom[88][10] = -32'd4198;
    weight_rom[88][11] = 32'd1566;
    weight_rom[88][12] = -32'd4255;
    weight_rom[88][13] = -32'd6394;
    weight_rom[88][14] = 32'd2475;
    weight_rom[88][15] = -32'd5696;
    weight_rom[88][16] = -32'd5512;
    weight_rom[88][17] = 32'd1403;
    weight_rom[88][18] = -32'd910;
    weight_rom[88][19] = 32'd2523;
    weight_rom[88][20] = -32'd881;
    weight_rom[88][21] = -32'd5978;
    weight_rom[88][22] = 32'd295;
    weight_rom[88][23] = 32'd3289;
    weight_rom[88][24] = -32'd735;
    weight_rom[88][25] = 32'd5266;
    weight_rom[88][26] = -32'd2453;
    weight_rom[88][27] = 32'd4779;
    weight_rom[88][28] = 32'd2943;
    weight_rom[88][29] = -32'd2669;
    weight_rom[88][30] = 32'd2464;
    weight_rom[88][31] = 32'd4173;
    weight_rom[88][32] = -32'd4807;
    weight_rom[88][33] = -32'd4923;
    weight_rom[88][34] = 32'd4906;
    weight_rom[88][35] = -32'd4743;
    weight_rom[88][36] = 32'd72;
    weight_rom[88][37] = 32'd583;
    weight_rom[88][38] = -32'd1286;
    weight_rom[88][39] = -32'd5571;
    weight_rom[88][40] = 32'd4843;
    weight_rom[88][41] = -32'd2164;
    weight_rom[88][42] = -32'd3056;
    weight_rom[88][43] = -32'd5687;
    weight_rom[88][44] = -32'd5181;
    weight_rom[88][45] = -32'd2359;
    weight_rom[88][46] = -32'd5900;
    weight_rom[88][47] = -32'd4893;
    weight_rom[88][48] = 32'd709;
    weight_rom[88][49] = -32'd5702;
    weight_rom[88][50] = -32'd991;
    weight_rom[88][51] = -32'd3936;
    weight_rom[88][52] = -32'd300;
    weight_rom[88][53] = 32'd1572;
    weight_rom[88][54] = -32'd6045;
    weight_rom[88][55] = -32'd2300;
    weight_rom[88][56] = -32'd5891;
    weight_rom[88][57] = 32'd2456;
    weight_rom[88][58] = -32'd6257;
    weight_rom[88][59] = -32'd655;
    weight_rom[88][60] = -32'd5204;
    weight_rom[88][61] = 32'd2700;
    weight_rom[88][62] = -32'd3537;
    weight_rom[88][63] = -32'd5201;
    weight_rom[89][0] = -32'd364;
    weight_rom[89][1] = 32'd3230;
    weight_rom[89][2] = 32'd1518;
    weight_rom[89][3] = 32'd5126;
    weight_rom[89][4] = -32'd2902;
    weight_rom[89][5] = -32'd4408;
    weight_rom[89][6] = -32'd366;
    weight_rom[89][7] = -32'd59;
    weight_rom[89][8] = 32'd484;
    weight_rom[89][9] = 32'd3625;
    weight_rom[89][10] = -32'd3440;
    weight_rom[89][11] = -32'd478;
    weight_rom[89][12] = 32'd2490;
    weight_rom[89][13] = -32'd3392;
    weight_rom[89][14] = 32'd4893;
    weight_rom[89][15] = -32'd162;
    weight_rom[89][16] = 32'd3034;
    weight_rom[89][17] = 32'd1721;
    weight_rom[89][18] = -32'd4684;
    weight_rom[89][19] = -32'd4791;
    weight_rom[89][20] = -32'd554;
    weight_rom[89][21] = -32'd4381;
    weight_rom[89][22] = -32'd5837;
    weight_rom[89][23] = -32'd5224;
    weight_rom[89][24] = -32'd6266;
    weight_rom[89][25] = -32'd3886;
    weight_rom[89][26] = 32'd2022;
    weight_rom[89][27] = -32'd4522;
    weight_rom[89][28] = -32'd5090;
    weight_rom[89][29] = 32'd5745;
    weight_rom[89][30] = -32'd4975;
    weight_rom[89][31] = -32'd6027;
    weight_rom[89][32] = 32'd1735;
    weight_rom[89][33] = 32'd4916;
    weight_rom[89][34] = 32'd4333;
    weight_rom[89][35] = 32'd4706;
    weight_rom[89][36] = 32'd101;
    weight_rom[89][37] = -32'd4458;
    weight_rom[89][38] = 32'd2277;
    weight_rom[89][39] = -32'd5162;
    weight_rom[89][40] = -32'd4185;
    weight_rom[89][41] = 32'd928;
    weight_rom[89][42] = 32'd77;
    weight_rom[89][43] = 32'd6194;
    weight_rom[89][44] = -32'd1009;
    weight_rom[89][45] = 32'd79;
    weight_rom[89][46] = -32'd4588;
    weight_rom[89][47] = -32'd4213;
    weight_rom[89][48] = -32'd4266;
    weight_rom[89][49] = -32'd449;
    weight_rom[89][50] = 32'd2814;
    weight_rom[89][51] = -32'd1687;
    weight_rom[89][52] = 32'd6482;
    weight_rom[89][53] = -32'd2094;
    weight_rom[89][54] = -32'd4105;
    weight_rom[89][55] = 32'd5834;
    weight_rom[89][56] = -32'd5978;
    weight_rom[89][57] = -32'd2288;
    weight_rom[89][58] = -32'd5074;
    weight_rom[89][59] = -32'd2192;
    weight_rom[89][60] = 32'd2870;
    weight_rom[89][61] = -32'd125;
    weight_rom[89][62] = -32'd1231;
    weight_rom[89][63] = 32'd5806;
    weight_rom[90][0] = -32'd4986;
    weight_rom[90][1] = 32'd1961;
    weight_rom[90][2] = 32'd1770;
    weight_rom[90][3] = 32'd363;
    weight_rom[90][4] = -32'd4233;
    weight_rom[90][5] = -32'd4400;
    weight_rom[90][6] = 32'd849;
    weight_rom[90][7] = 32'd2469;
    weight_rom[90][8] = 32'd1218;
    weight_rom[90][9] = 32'd3551;
    weight_rom[90][10] = 32'd6178;
    weight_rom[90][11] = -32'd1575;
    weight_rom[90][12] = -32'd3919;
    weight_rom[90][13] = 32'd6237;
    weight_rom[90][14] = 32'd1786;
    weight_rom[90][15] = -32'd6113;
    weight_rom[90][16] = -32'd4097;
    weight_rom[90][17] = 32'd1201;
    weight_rom[90][18] = 32'd5113;
    weight_rom[90][19] = -32'd2629;
    weight_rom[90][20] = -32'd3815;
    weight_rom[90][21] = -32'd713;
    weight_rom[90][22] = 32'd6200;
    weight_rom[90][23] = -32'd2911;
    weight_rom[90][24] = -32'd2607;
    weight_rom[90][25] = -32'd5675;
    weight_rom[90][26] = -32'd3512;
    weight_rom[90][27] = -32'd5469;
    weight_rom[90][28] = 32'd1419;
    weight_rom[90][29] = 32'd4177;
    weight_rom[90][30] = 32'd5747;
    weight_rom[90][31] = 32'd5110;
    weight_rom[90][32] = -32'd4871;
    weight_rom[90][33] = 32'd6172;
    weight_rom[90][34] = -32'd3609;
    weight_rom[90][35] = 32'd0;
    weight_rom[90][36] = -32'd4739;
    weight_rom[90][37] = 32'd2506;
    weight_rom[90][38] = -32'd650;
    weight_rom[90][39] = 32'd4423;
    weight_rom[90][40] = 32'd5867;
    weight_rom[90][41] = 32'd5368;
    weight_rom[90][42] = 32'd3640;
    weight_rom[90][43] = -32'd1834;
    weight_rom[90][44] = 32'd3874;
    weight_rom[90][45] = -32'd4423;
    weight_rom[90][46] = 32'd492;
    weight_rom[90][47] = -32'd91;
    weight_rom[90][48] = -32'd1589;
    weight_rom[90][49] = -32'd3404;
    weight_rom[90][50] = 32'd1360;
    weight_rom[90][51] = 32'd22;
    weight_rom[90][52] = 32'd2348;
    weight_rom[90][53] = 32'd4665;
    weight_rom[90][54] = 32'd4341;
    weight_rom[90][55] = -32'd2848;
    weight_rom[90][56] = 32'd2888;
    weight_rom[90][57] = -32'd5311;
    weight_rom[90][58] = 32'd1434;
    weight_rom[90][59] = -32'd808;
    weight_rom[90][60] = 32'd50;
    weight_rom[90][61] = -32'd3175;
    weight_rom[90][62] = 32'd4275;
    weight_rom[90][63] = 32'd3867;
    weight_rom[91][0] = 32'd2795;
    weight_rom[91][1] = 32'd4577;
    weight_rom[91][2] = -32'd5959;
    weight_rom[91][3] = 32'd6461;
    weight_rom[91][4] = -32'd5390;
    weight_rom[91][5] = 32'd4123;
    weight_rom[91][6] = -32'd5692;
    weight_rom[91][7] = -32'd854;
    weight_rom[91][8] = 32'd1049;
    weight_rom[91][9] = 32'd4519;
    weight_rom[91][10] = -32'd4181;
    weight_rom[91][11] = 32'd4762;
    weight_rom[91][12] = 32'd469;
    weight_rom[91][13] = 32'd3952;
    weight_rom[91][14] = 32'd3422;
    weight_rom[91][15] = -32'd5732;
    weight_rom[91][16] = 32'd4694;
    weight_rom[91][17] = 32'd2655;
    weight_rom[91][18] = -32'd2020;
    weight_rom[91][19] = -32'd1851;
    weight_rom[91][20] = -32'd1720;
    weight_rom[91][21] = -32'd3811;
    weight_rom[91][22] = -32'd3589;
    weight_rom[91][23] = -32'd2931;
    weight_rom[91][24] = 32'd34;
    weight_rom[91][25] = 32'd4946;
    weight_rom[91][26] = -32'd6365;
    weight_rom[91][27] = -32'd202;
    weight_rom[91][28] = -32'd2869;
    weight_rom[91][29] = 32'd6338;
    weight_rom[91][30] = -32'd4178;
    weight_rom[91][31] = 32'd6448;
    weight_rom[91][32] = 32'd1028;
    weight_rom[91][33] = -32'd4231;
    weight_rom[91][34] = -32'd1319;
    weight_rom[91][35] = 32'd2292;
    weight_rom[91][36] = 32'd6327;
    weight_rom[91][37] = -32'd4357;
    weight_rom[91][38] = 32'd3263;
    weight_rom[91][39] = -32'd3410;
    weight_rom[91][40] = -32'd3686;
    weight_rom[91][41] = -32'd6472;
    weight_rom[91][42] = 32'd4696;
    weight_rom[91][43] = -32'd290;
    weight_rom[91][44] = -32'd4700;
    weight_rom[91][45] = 32'd6025;
    weight_rom[91][46] = 32'd993;
    weight_rom[91][47] = -32'd5479;
    weight_rom[91][48] = 32'd4497;
    weight_rom[91][49] = -32'd395;
    weight_rom[91][50] = -32'd2635;
    weight_rom[91][51] = 32'd2955;
    weight_rom[91][52] = -32'd5582;
    weight_rom[91][53] = -32'd856;
    weight_rom[91][54] = 32'd3496;
    weight_rom[91][55] = -32'd512;
    weight_rom[91][56] = -32'd727;
    weight_rom[91][57] = 32'd6237;
    weight_rom[91][58] = 32'd4201;
    weight_rom[91][59] = -32'd3110;
    weight_rom[91][60] = 32'd2736;
    weight_rom[91][61] = 32'd5045;
    weight_rom[91][62] = -32'd3569;
    weight_rom[91][63] = -32'd4177;
    weight_rom[92][0] = 32'd3418;
    weight_rom[92][1] = 32'd2065;
    weight_rom[92][2] = -32'd1643;
    weight_rom[92][3] = -32'd5586;
    weight_rom[92][4] = -32'd4972;
    weight_rom[92][5] = 32'd2165;
    weight_rom[92][6] = 32'd3611;
    weight_rom[92][7] = -32'd3323;
    weight_rom[92][8] = -32'd5354;
    weight_rom[92][9] = 32'd3421;
    weight_rom[92][10] = 32'd4644;
    weight_rom[92][11] = 32'd250;
    weight_rom[92][12] = -32'd5286;
    weight_rom[92][13] = 32'd6023;
    weight_rom[92][14] = -32'd4455;
    weight_rom[92][15] = 32'd5327;
    weight_rom[92][16] = 32'd4182;
    weight_rom[92][17] = -32'd3441;
    weight_rom[92][18] = -32'd4529;
    weight_rom[92][19] = 32'd3990;
    weight_rom[92][20] = -32'd1706;
    weight_rom[92][21] = -32'd5898;
    weight_rom[92][22] = -32'd2566;
    weight_rom[92][23] = -32'd891;
    weight_rom[92][24] = -32'd5817;
    weight_rom[92][25] = -32'd1449;
    weight_rom[92][26] = 32'd3464;
    weight_rom[92][27] = -32'd2589;
    weight_rom[92][28] = -32'd4279;
    weight_rom[92][29] = -32'd3150;
    weight_rom[92][30] = 32'd1608;
    weight_rom[92][31] = -32'd2699;
    weight_rom[92][32] = 32'd2535;
    weight_rom[92][33] = 32'd2910;
    weight_rom[92][34] = -32'd1183;
    weight_rom[92][35] = -32'd3420;
    weight_rom[92][36] = -32'd3277;
    weight_rom[92][37] = -32'd2486;
    weight_rom[92][38] = -32'd1874;
    weight_rom[92][39] = -32'd3998;
    weight_rom[92][40] = -32'd2277;
    weight_rom[92][41] = 32'd4072;
    weight_rom[92][42] = 32'd4520;
    weight_rom[92][43] = -32'd1896;
    weight_rom[92][44] = -32'd4845;
    weight_rom[92][45] = 32'd4608;
    weight_rom[92][46] = 32'd1902;
    weight_rom[92][47] = -32'd3984;
    weight_rom[92][48] = 32'd1890;
    weight_rom[92][49] = -32'd583;
    weight_rom[92][50] = -32'd1168;
    weight_rom[92][51] = -32'd5069;
    weight_rom[92][52] = 32'd6459;
    weight_rom[92][53] = -32'd4026;
    weight_rom[92][54] = -32'd1957;
    weight_rom[92][55] = 32'd2245;
    weight_rom[92][56] = -32'd3194;
    weight_rom[92][57] = -32'd2801;
    weight_rom[92][58] = -32'd2814;
    weight_rom[92][59] = -32'd4394;
    weight_rom[92][60] = -32'd3290;
    weight_rom[92][61] = 32'd1009;
    weight_rom[92][62] = 32'd320;
    weight_rom[92][63] = 32'd2778;
    weight_rom[93][0] = 32'd803;
    weight_rom[93][1] = 32'd895;
    weight_rom[93][2] = 32'd1649;
    weight_rom[93][3] = 32'd705;
    weight_rom[93][4] = -32'd514;
    weight_rom[93][5] = 32'd302;
    weight_rom[93][6] = -32'd612;
    weight_rom[93][7] = 32'd4182;
    weight_rom[93][8] = 32'd4947;
    weight_rom[93][9] = 32'd1654;
    weight_rom[93][10] = -32'd101;
    weight_rom[93][11] = -32'd272;
    weight_rom[93][12] = -32'd650;
    weight_rom[93][13] = -32'd159;
    weight_rom[93][14] = -32'd503;
    weight_rom[93][15] = -32'd4728;
    weight_rom[93][16] = 32'd534;
    weight_rom[93][17] = 32'd162;
    weight_rom[93][18] = -32'd6220;
    weight_rom[93][19] = -32'd2899;
    weight_rom[93][20] = -32'd5867;
    weight_rom[93][21] = 32'd4504;
    weight_rom[93][22] = -32'd2569;
    weight_rom[93][23] = 32'd6296;
    weight_rom[93][24] = -32'd116;
    weight_rom[93][25] = 32'd547;
    weight_rom[93][26] = 32'd1621;
    weight_rom[93][27] = 32'd831;
    weight_rom[93][28] = -32'd1576;
    weight_rom[93][29] = 32'd6156;
    weight_rom[93][30] = -32'd3634;
    weight_rom[93][31] = -32'd3796;
    weight_rom[93][32] = 32'd2629;
    weight_rom[93][33] = -32'd6025;
    weight_rom[93][34] = 32'd6268;
    weight_rom[93][35] = 32'd3382;
    weight_rom[93][36] = -32'd5591;
    weight_rom[93][37] = 32'd43;
    weight_rom[93][38] = 32'd1766;
    weight_rom[93][39] = 32'd64;
    weight_rom[93][40] = 32'd3357;
    weight_rom[93][41] = 32'd5876;
    weight_rom[93][42] = -32'd1839;
    weight_rom[93][43] = 32'd2392;
    weight_rom[93][44] = 32'd1879;
    weight_rom[93][45] = 32'd4768;
    weight_rom[93][46] = -32'd6331;
    weight_rom[93][47] = 32'd5816;
    weight_rom[93][48] = 32'd1975;
    weight_rom[93][49] = 32'd1076;
    weight_rom[93][50] = -32'd3700;
    weight_rom[93][51] = -32'd1227;
    weight_rom[93][52] = -32'd1207;
    weight_rom[93][53] = -32'd4048;
    weight_rom[93][54] = -32'd1614;
    weight_rom[93][55] = -32'd4427;
    weight_rom[93][56] = -32'd4057;
    weight_rom[93][57] = -32'd998;
    weight_rom[93][58] = -32'd3418;
    weight_rom[93][59] = 32'd2479;
    weight_rom[93][60] = -32'd2301;
    weight_rom[93][61] = -32'd3654;
    weight_rom[93][62] = 32'd4012;
    weight_rom[93][63] = -32'd1507;
    weight_rom[94][0] = 32'd3551;
    weight_rom[94][1] = -32'd5325;
    weight_rom[94][2] = 32'd41;
    weight_rom[94][3] = 32'd6151;
    weight_rom[94][4] = -32'd3849;
    weight_rom[94][5] = -32'd1850;
    weight_rom[94][6] = 32'd319;
    weight_rom[94][7] = 32'd3924;
    weight_rom[94][8] = -32'd3072;
    weight_rom[94][9] = -32'd4833;
    weight_rom[94][10] = -32'd3313;
    weight_rom[94][11] = -32'd6217;
    weight_rom[94][12] = 32'd3357;
    weight_rom[94][13] = -32'd5115;
    weight_rom[94][14] = -32'd6431;
    weight_rom[94][15] = 32'd424;
    weight_rom[94][16] = 32'd2755;
    weight_rom[94][17] = -32'd5187;
    weight_rom[94][18] = 32'd1911;
    weight_rom[94][19] = -32'd3791;
    weight_rom[94][20] = 32'd3507;
    weight_rom[94][21] = 32'd6307;
    weight_rom[94][22] = -32'd3533;
    weight_rom[94][23] = -32'd5668;
    weight_rom[94][24] = 32'd5598;
    weight_rom[94][25] = 32'd6135;
    weight_rom[94][26] = 32'd3438;
    weight_rom[94][27] = 32'd3982;
    weight_rom[94][28] = 32'd3951;
    weight_rom[94][29] = -32'd901;
    weight_rom[94][30] = -32'd2526;
    weight_rom[94][31] = 32'd3478;
    weight_rom[94][32] = 32'd3322;
    weight_rom[94][33] = -32'd1239;
    weight_rom[94][34] = -32'd4182;
    weight_rom[94][35] = 32'd3407;
    weight_rom[94][36] = 32'd2138;
    weight_rom[94][37] = 32'd3885;
    weight_rom[94][38] = -32'd4110;
    weight_rom[94][39] = 32'd3522;
    weight_rom[94][40] = -32'd1392;
    weight_rom[94][41] = -32'd5356;
    weight_rom[94][42] = 32'd2454;
    weight_rom[94][43] = 32'd2126;
    weight_rom[94][44] = -32'd3969;
    weight_rom[94][45] = -32'd1221;
    weight_rom[94][46] = 32'd6034;
    weight_rom[94][47] = 32'd6245;
    weight_rom[94][48] = 32'd4807;
    weight_rom[94][49] = -32'd1877;
    weight_rom[94][50] = 32'd6108;
    weight_rom[94][51] = -32'd195;
    weight_rom[94][52] = -32'd2786;
    weight_rom[94][53] = 32'd3522;
    weight_rom[94][54] = 32'd439;
    weight_rom[94][55] = -32'd177;
    weight_rom[94][56] = 32'd2227;
    weight_rom[94][57] = 32'd1964;
    weight_rom[94][58] = 32'd3761;
    weight_rom[94][59] = 32'd190;
    weight_rom[94][60] = -32'd2172;
    weight_rom[94][61] = -32'd3026;
    weight_rom[94][62] = -32'd1920;
    weight_rom[94][63] = -32'd1280;
    weight_rom[95][0] = -32'd81;
    weight_rom[95][1] = -32'd1733;
    weight_rom[95][2] = 32'd4672;
    weight_rom[95][3] = 32'd302;
    weight_rom[95][4] = -32'd1779;
    weight_rom[95][5] = 32'd4944;
    weight_rom[95][6] = -32'd776;
    weight_rom[95][7] = 32'd2551;
    weight_rom[95][8] = -32'd4856;
    weight_rom[95][9] = -32'd6127;
    weight_rom[95][10] = 32'd4859;
    weight_rom[95][11] = -32'd2080;
    weight_rom[95][12] = -32'd1997;
    weight_rom[95][13] = 32'd628;
    weight_rom[95][14] = -32'd3320;
    weight_rom[95][15] = -32'd1165;
    weight_rom[95][16] = -32'd2433;
    weight_rom[95][17] = -32'd1513;
    weight_rom[95][18] = 32'd1794;
    weight_rom[95][19] = 32'd5995;
    weight_rom[95][20] = -32'd1094;
    weight_rom[95][21] = 32'd3842;
    weight_rom[95][22] = -32'd6534;
    weight_rom[95][23] = 32'd245;
    weight_rom[95][24] = -32'd5172;
    weight_rom[95][25] = -32'd5681;
    weight_rom[95][26] = -32'd6043;
    weight_rom[95][27] = -32'd4755;
    weight_rom[95][28] = -32'd1414;
    weight_rom[95][29] = -32'd1998;
    weight_rom[95][30] = 32'd608;
    weight_rom[95][31] = -32'd3237;
    weight_rom[95][32] = 32'd4887;
    weight_rom[95][33] = 32'd213;
    weight_rom[95][34] = 32'd3921;
    weight_rom[95][35] = -32'd2456;
    weight_rom[95][36] = 32'd1249;
    weight_rom[95][37] = 32'd3138;
    weight_rom[95][38] = 32'd3268;
    weight_rom[95][39] = -32'd5741;
    weight_rom[95][40] = 32'd1418;
    weight_rom[95][41] = -32'd4437;
    weight_rom[95][42] = -32'd2453;
    weight_rom[95][43] = 32'd2822;
    weight_rom[95][44] = -32'd5274;
    weight_rom[95][45] = 32'd3438;
    weight_rom[95][46] = -32'd5969;
    weight_rom[95][47] = -32'd1621;
    weight_rom[95][48] = 32'd5163;
    weight_rom[95][49] = -32'd4400;
    weight_rom[95][50] = -32'd4841;
    weight_rom[95][51] = 32'd535;
    weight_rom[95][52] = 32'd758;
    weight_rom[95][53] = -32'd3072;
    weight_rom[95][54] = -32'd6550;
    weight_rom[95][55] = 32'd3126;
    weight_rom[95][56] = -32'd6548;
    weight_rom[95][57] = -32'd6229;
    weight_rom[95][58] = -32'd5814;
    weight_rom[95][59] = -32'd3930;
    weight_rom[95][60] = -32'd6216;
    weight_rom[95][61] = 32'd3973;
    weight_rom[95][62] = 32'd1863;
    weight_rom[95][63] = 32'd3713;
    weight_rom[96][0] = 32'd297;
    weight_rom[96][1] = -32'd3077;
    weight_rom[96][2] = 32'd2080;
    weight_rom[96][3] = 32'd1696;
    weight_rom[96][4] = 32'd44;
    weight_rom[96][5] = -32'd1409;
    weight_rom[96][6] = -32'd1300;
    weight_rom[96][7] = -32'd2986;
    weight_rom[96][8] = 32'd5095;
    weight_rom[96][9] = 32'd5516;
    weight_rom[96][10] = -32'd716;
    weight_rom[96][11] = -32'd1570;
    weight_rom[96][12] = 32'd2161;
    weight_rom[96][13] = -32'd598;
    weight_rom[96][14] = 32'd2968;
    weight_rom[96][15] = -32'd2000;
    weight_rom[96][16] = -32'd377;
    weight_rom[96][17] = -32'd161;
    weight_rom[96][18] = -32'd2089;
    weight_rom[96][19] = -32'd6437;
    weight_rom[96][20] = 32'd4222;
    weight_rom[96][21] = 32'd4637;
    weight_rom[96][22] = 32'd3006;
    weight_rom[96][23] = -32'd4202;
    weight_rom[96][24] = 32'd3466;
    weight_rom[96][25] = 32'd1944;
    weight_rom[96][26] = 32'd4418;
    weight_rom[96][27] = 32'd1057;
    weight_rom[96][28] = 32'd3286;
    weight_rom[96][29] = -32'd5893;
    weight_rom[96][30] = -32'd1085;
    weight_rom[96][31] = 32'd4791;
    weight_rom[96][32] = 32'd0;
    weight_rom[96][33] = 32'd1057;
    weight_rom[96][34] = -32'd2173;
    weight_rom[96][35] = -32'd1170;
    weight_rom[96][36] = -32'd1112;
    weight_rom[96][37] = 32'd1907;
    weight_rom[96][38] = 32'd598;
    weight_rom[96][39] = 32'd1006;
    weight_rom[96][40] = -32'd726;
    weight_rom[96][41] = 32'd6039;
    weight_rom[96][42] = -32'd5755;
    weight_rom[96][43] = -32'd3038;
    weight_rom[96][44] = -32'd4366;
    weight_rom[96][45] = -32'd4667;
    weight_rom[96][46] = -32'd4678;
    weight_rom[96][47] = 32'd5548;
    weight_rom[96][48] = 32'd5502;
    weight_rom[96][49] = 32'd48;
    weight_rom[96][50] = -32'd1679;
    weight_rom[96][51] = 32'd4172;
    weight_rom[96][52] = -32'd2564;
    weight_rom[96][53] = 32'd3502;
    weight_rom[96][54] = -32'd3391;
    weight_rom[96][55] = 32'd4808;
    weight_rom[96][56] = 32'd4009;
    weight_rom[96][57] = 32'd4066;
    weight_rom[96][58] = -32'd1711;
    weight_rom[96][59] = -32'd2364;
    weight_rom[96][60] = -32'd2083;
    weight_rom[96][61] = -32'd5974;
    weight_rom[96][62] = -32'd3334;
    weight_rom[96][63] = 32'd6065;
    weight_rom[97][0] = -32'd949;
    weight_rom[97][1] = -32'd3355;
    weight_rom[97][2] = -32'd4417;
    weight_rom[97][3] = 32'd2565;
    weight_rom[97][4] = 32'd2495;
    weight_rom[97][5] = 32'd4149;
    weight_rom[97][6] = 32'd781;
    weight_rom[97][7] = 32'd1182;
    weight_rom[97][8] = 32'd5972;
    weight_rom[97][9] = 32'd1528;
    weight_rom[97][10] = 32'd194;
    weight_rom[97][11] = -32'd1326;
    weight_rom[97][12] = 32'd3872;
    weight_rom[97][13] = 32'd4513;
    weight_rom[97][14] = 32'd6446;
    weight_rom[97][15] = 32'd5240;
    weight_rom[97][16] = 32'd4215;
    weight_rom[97][17] = 32'd1995;
    weight_rom[97][18] = -32'd5613;
    weight_rom[97][19] = 32'd6525;
    weight_rom[97][20] = 32'd4592;
    weight_rom[97][21] = -32'd3381;
    weight_rom[97][22] = 32'd6119;
    weight_rom[97][23] = 32'd6169;
    weight_rom[97][24] = -32'd1183;
    weight_rom[97][25] = -32'd5582;
    weight_rom[97][26] = 32'd1566;
    weight_rom[97][27] = 32'd72;
    weight_rom[97][28] = -32'd4908;
    weight_rom[97][29] = -32'd5861;
    weight_rom[97][30] = -32'd4453;
    weight_rom[97][31] = -32'd5205;
    weight_rom[97][32] = 32'd3017;
    weight_rom[97][33] = 32'd5713;
    weight_rom[97][34] = 32'd3026;
    weight_rom[97][35] = -32'd3805;
    weight_rom[97][36] = -32'd1019;
    weight_rom[97][37] = -32'd4511;
    weight_rom[97][38] = -32'd3878;
    weight_rom[97][39] = -32'd4991;
    weight_rom[97][40] = 32'd3176;
    weight_rom[97][41] = 32'd492;
    weight_rom[97][42] = 32'd2641;
    weight_rom[97][43] = -32'd2416;
    weight_rom[97][44] = 32'd5553;
    weight_rom[97][45] = -32'd6440;
    weight_rom[97][46] = -32'd6369;
    weight_rom[97][47] = 32'd587;
    weight_rom[97][48] = -32'd5310;
    weight_rom[97][49] = 32'd4328;
    weight_rom[97][50] = -32'd6214;
    weight_rom[97][51] = -32'd4303;
    weight_rom[97][52] = -32'd5420;
    weight_rom[97][53] = -32'd3855;
    weight_rom[97][54] = -32'd3824;
    weight_rom[97][55] = 32'd1654;
    weight_rom[97][56] = -32'd5514;
    weight_rom[97][57] = 32'd479;
    weight_rom[97][58] = 32'd76;
    weight_rom[97][59] = 32'd1203;
    weight_rom[97][60] = 32'd3975;
    weight_rom[97][61] = 32'd6449;
    weight_rom[97][62] = -32'd5121;
    weight_rom[97][63] = -32'd4893;
    weight_rom[98][0] = -32'd6220;
    weight_rom[98][1] = 32'd6199;
    weight_rom[98][2] = -32'd5628;
    weight_rom[98][3] = -32'd595;
    weight_rom[98][4] = -32'd6038;
    weight_rom[98][5] = -32'd797;
    weight_rom[98][6] = -32'd4518;
    weight_rom[98][7] = -32'd1822;
    weight_rom[98][8] = 32'd4746;
    weight_rom[98][9] = 32'd3886;
    weight_rom[98][10] = -32'd1845;
    weight_rom[98][11] = 32'd1050;
    weight_rom[98][12] = 32'd5599;
    weight_rom[98][13] = -32'd5267;
    weight_rom[98][14] = -32'd5253;
    weight_rom[98][15] = -32'd6267;
    weight_rom[98][16] = -32'd533;
    weight_rom[98][17] = 32'd5905;
    weight_rom[98][18] = -32'd1184;
    weight_rom[98][19] = 32'd2317;
    weight_rom[98][20] = -32'd3774;
    weight_rom[98][21] = 32'd6037;
    weight_rom[98][22] = -32'd3613;
    weight_rom[98][23] = -32'd5068;
    weight_rom[98][24] = 32'd2033;
    weight_rom[98][25] = -32'd1632;
    weight_rom[98][26] = 32'd830;
    weight_rom[98][27] = -32'd4665;
    weight_rom[98][28] = 32'd3575;
    weight_rom[98][29] = 32'd2516;
    weight_rom[98][30] = -32'd4313;
    weight_rom[98][31] = -32'd4902;
    weight_rom[98][32] = 32'd1562;
    weight_rom[98][33] = 32'd2257;
    weight_rom[98][34] = -32'd1048;
    weight_rom[98][35] = 32'd6246;
    weight_rom[98][36] = 32'd3736;
    weight_rom[98][37] = 32'd616;
    weight_rom[98][38] = -32'd2727;
    weight_rom[98][39] = -32'd6075;
    weight_rom[98][40] = -32'd3560;
    weight_rom[98][41] = -32'd6367;
    weight_rom[98][42] = -32'd6424;
    weight_rom[98][43] = -32'd4911;
    weight_rom[98][44] = 32'd4213;
    weight_rom[98][45] = -32'd6291;
    weight_rom[98][46] = 32'd876;
    weight_rom[98][47] = -32'd3018;
    weight_rom[98][48] = 32'd578;
    weight_rom[98][49] = 32'd2149;
    weight_rom[98][50] = -32'd3646;
    weight_rom[98][51] = 32'd4034;
    weight_rom[98][52] = -32'd6534;
    weight_rom[98][53] = -32'd2337;
    weight_rom[98][54] = -32'd3270;
    weight_rom[98][55] = 32'd2215;
    weight_rom[98][56] = -32'd4043;
    weight_rom[98][57] = -32'd2906;
    weight_rom[98][58] = 32'd791;
    weight_rom[98][59] = -32'd5606;
    weight_rom[98][60] = 32'd5207;
    weight_rom[98][61] = -32'd4845;
    weight_rom[98][62] = 32'd3858;
    weight_rom[98][63] = -32'd1040;
    weight_rom[99][0] = -32'd5139;
    weight_rom[99][1] = -32'd1401;
    weight_rom[99][2] = 32'd1866;
    weight_rom[99][3] = 32'd1671;
    weight_rom[99][4] = 32'd3924;
    weight_rom[99][5] = -32'd1612;
    weight_rom[99][6] = -32'd4169;
    weight_rom[99][7] = -32'd5353;
    weight_rom[99][8] = 32'd4056;
    weight_rom[99][9] = -32'd242;
    weight_rom[99][10] = 32'd1218;
    weight_rom[99][11] = 32'd440;
    weight_rom[99][12] = -32'd3478;
    weight_rom[99][13] = -32'd154;
    weight_rom[99][14] = -32'd1291;
    weight_rom[99][15] = 32'd2146;
    weight_rom[99][16] = -32'd1863;
    weight_rom[99][17] = 32'd1319;
    weight_rom[99][18] = -32'd2474;
    weight_rom[99][19] = 32'd4305;
    weight_rom[99][20] = 32'd2062;
    weight_rom[99][21] = -32'd3972;
    weight_rom[99][22] = 32'd2137;
    weight_rom[99][23] = -32'd1263;
    weight_rom[99][24] = -32'd3142;
    weight_rom[99][25] = 32'd3982;
    weight_rom[99][26] = 32'd1633;
    weight_rom[99][27] = 32'd1625;
    weight_rom[99][28] = -32'd3448;
    weight_rom[99][29] = -32'd551;
    weight_rom[99][30] = -32'd1072;
    weight_rom[99][31] = 32'd6280;
    weight_rom[99][32] = -32'd4107;
    weight_rom[99][33] = -32'd245;
    weight_rom[99][34] = 32'd1027;
    weight_rom[99][35] = 32'd1908;
    weight_rom[99][36] = -32'd3988;
    weight_rom[99][37] = -32'd5407;
    weight_rom[99][38] = 32'd3258;
    weight_rom[99][39] = -32'd5862;
    weight_rom[99][40] = -32'd5787;
    weight_rom[99][41] = -32'd3176;
    weight_rom[99][42] = -32'd1190;
    weight_rom[99][43] = 32'd2038;
    weight_rom[99][44] = -32'd1912;
    weight_rom[99][45] = 32'd1135;
    weight_rom[99][46] = 32'd5665;
    weight_rom[99][47] = 32'd2652;
    weight_rom[99][48] = 32'd3152;
    weight_rom[99][49] = -32'd2118;
    weight_rom[99][50] = 32'd3676;
    weight_rom[99][51] = 32'd2528;
    weight_rom[99][52] = -32'd660;
    weight_rom[99][53] = -32'd452;
    weight_rom[99][54] = 32'd4009;
    weight_rom[99][55] = -32'd4898;
    weight_rom[99][56] = -32'd1491;
    weight_rom[99][57] = -32'd5746;
    weight_rom[99][58] = 32'd2996;
    weight_rom[99][59] = -32'd4620;
    weight_rom[99][60] = 32'd238;
    weight_rom[99][61] = 32'd3880;
    weight_rom[99][62] = -32'd5256;
    weight_rom[99][63] = -32'd249;
    weight_rom[100][0] = -32'd6141;
    weight_rom[100][1] = 32'd5138;
    weight_rom[100][2] = -32'd6206;
    weight_rom[100][3] = 32'd1105;
    weight_rom[100][4] = 32'd1676;
    weight_rom[100][5] = -32'd489;
    weight_rom[100][6] = 32'd4741;
    weight_rom[100][7] = 32'd5469;
    weight_rom[100][8] = 32'd2034;
    weight_rom[100][9] = -32'd5015;
    weight_rom[100][10] = -32'd4410;
    weight_rom[100][11] = 32'd1414;
    weight_rom[100][12] = -32'd1319;
    weight_rom[100][13] = -32'd4586;
    weight_rom[100][14] = 32'd3933;
    weight_rom[100][15] = 32'd6073;
    weight_rom[100][16] = -32'd75;
    weight_rom[100][17] = 32'd3192;
    weight_rom[100][18] = 32'd2321;
    weight_rom[100][19] = -32'd2691;
    weight_rom[100][20] = -32'd363;
    weight_rom[100][21] = 32'd5916;
    weight_rom[100][22] = 32'd3170;
    weight_rom[100][23] = 32'd3118;
    weight_rom[100][24] = -32'd4463;
    weight_rom[100][25] = -32'd872;
    weight_rom[100][26] = 32'd4776;
    weight_rom[100][27] = -32'd2966;
    weight_rom[100][28] = 32'd2325;
    weight_rom[100][29] = -32'd3584;
    weight_rom[100][30] = 32'd3372;
    weight_rom[100][31] = 32'd2278;
    weight_rom[100][32] = -32'd6216;
    weight_rom[100][33] = 32'd4058;
    weight_rom[100][34] = 32'd4359;
    weight_rom[100][35] = 32'd5695;
    weight_rom[100][36] = 32'd4197;
    weight_rom[100][37] = -32'd1607;
    weight_rom[100][38] = -32'd228;
    weight_rom[100][39] = 32'd4379;
    weight_rom[100][40] = -32'd2622;
    weight_rom[100][41] = -32'd656;
    weight_rom[100][42] = -32'd2236;
    weight_rom[100][43] = -32'd6031;
    weight_rom[100][44] = 32'd2042;
    weight_rom[100][45] = -32'd584;
    weight_rom[100][46] = 32'd2175;
    weight_rom[100][47] = 32'd2082;
    weight_rom[100][48] = 32'd3367;
    weight_rom[100][49] = 32'd5708;
    weight_rom[100][50] = -32'd3916;
    weight_rom[100][51] = 32'd732;
    weight_rom[100][52] = 32'd4415;
    weight_rom[100][53] = 32'd5809;
    weight_rom[100][54] = -32'd2887;
    weight_rom[100][55] = 32'd5842;
    weight_rom[100][56] = -32'd198;
    weight_rom[100][57] = -32'd4423;
    weight_rom[100][58] = -32'd1902;
    weight_rom[100][59] = -32'd5593;
    weight_rom[100][60] = -32'd583;
    weight_rom[100][61] = -32'd1379;
    weight_rom[100][62] = -32'd2996;
    weight_rom[100][63] = -32'd1621;
    weight_rom[101][0] = 32'd1787;
    weight_rom[101][1] = 32'd1718;
    weight_rom[101][2] = 32'd1124;
    weight_rom[101][3] = 32'd5258;
    weight_rom[101][4] = -32'd5481;
    weight_rom[101][5] = -32'd2603;
    weight_rom[101][6] = 32'd5847;
    weight_rom[101][7] = -32'd4760;
    weight_rom[101][8] = 32'd666;
    weight_rom[101][9] = -32'd4912;
    weight_rom[101][10] = -32'd1427;
    weight_rom[101][11] = 32'd3471;
    weight_rom[101][12] = -32'd4555;
    weight_rom[101][13] = -32'd2298;
    weight_rom[101][14] = -32'd3879;
    weight_rom[101][15] = 32'd788;
    weight_rom[101][16] = 32'd4302;
    weight_rom[101][17] = 32'd82;
    weight_rom[101][18] = 32'd1386;
    weight_rom[101][19] = -32'd6365;
    weight_rom[101][20] = 32'd4982;
    weight_rom[101][21] = 32'd6485;
    weight_rom[101][22] = 32'd4566;
    weight_rom[101][23] = 32'd2681;
    weight_rom[101][24] = -32'd4450;
    weight_rom[101][25] = 32'd6516;
    weight_rom[101][26] = 32'd1139;
    weight_rom[101][27] = -32'd159;
    weight_rom[101][28] = 32'd862;
    weight_rom[101][29] = 32'd1493;
    weight_rom[101][30] = 32'd5216;
    weight_rom[101][31] = 32'd4546;
    weight_rom[101][32] = -32'd2824;
    weight_rom[101][33] = 32'd5905;
    weight_rom[101][34] = 32'd3986;
    weight_rom[101][35] = -32'd2577;
    weight_rom[101][36] = 32'd1949;
    weight_rom[101][37] = -32'd1133;
    weight_rom[101][38] = -32'd3722;
    weight_rom[101][39] = -32'd5007;
    weight_rom[101][40] = -32'd336;
    weight_rom[101][41] = 32'd2528;
    weight_rom[101][42] = 32'd2534;
    weight_rom[101][43] = 32'd1280;
    weight_rom[101][44] = 32'd488;
    weight_rom[101][45] = 32'd236;
    weight_rom[101][46] = 32'd4229;
    weight_rom[101][47] = 32'd6411;
    weight_rom[101][48] = 32'd1398;
    weight_rom[101][49] = 32'd5402;
    weight_rom[101][50] = -32'd5504;
    weight_rom[101][51] = 32'd2615;
    weight_rom[101][52] = 32'd947;
    weight_rom[101][53] = 32'd5658;
    weight_rom[101][54] = -32'd4043;
    weight_rom[101][55] = -32'd4815;
    weight_rom[101][56] = -32'd1900;
    weight_rom[101][57] = 32'd5177;
    weight_rom[101][58] = 32'd1476;
    weight_rom[101][59] = 32'd4093;
    weight_rom[101][60] = -32'd6149;
    weight_rom[101][61] = -32'd102;
    weight_rom[101][62] = 32'd4654;
    weight_rom[101][63] = -32'd1793;
    weight_rom[102][0] = -32'd2433;
    weight_rom[102][1] = 32'd3864;
    weight_rom[102][2] = 32'd5770;
    weight_rom[102][3] = -32'd5957;
    weight_rom[102][4] = 32'd4896;
    weight_rom[102][5] = 32'd3245;
    weight_rom[102][6] = -32'd1660;
    weight_rom[102][7] = 32'd5901;
    weight_rom[102][8] = -32'd5413;
    weight_rom[102][9] = 32'd2432;
    weight_rom[102][10] = 32'd6152;
    weight_rom[102][11] = 32'd4102;
    weight_rom[102][12] = 32'd6455;
    weight_rom[102][13] = 32'd3111;
    weight_rom[102][14] = 32'd722;
    weight_rom[102][15] = 32'd5725;
    weight_rom[102][16] = -32'd2159;
    weight_rom[102][17] = 32'd1757;
    weight_rom[102][18] = -32'd1774;
    weight_rom[102][19] = 32'd3117;
    weight_rom[102][20] = -32'd3725;
    weight_rom[102][21] = 32'd2775;
    weight_rom[102][22] = -32'd1014;
    weight_rom[102][23] = -32'd1012;
    weight_rom[102][24] = -32'd5629;
    weight_rom[102][25] = 32'd774;
    weight_rom[102][26] = 32'd1061;
    weight_rom[102][27] = -32'd5475;
    weight_rom[102][28] = 32'd5624;
    weight_rom[102][29] = -32'd3239;
    weight_rom[102][30] = -32'd5450;
    weight_rom[102][31] = -32'd2302;
    weight_rom[102][32] = -32'd746;
    weight_rom[102][33] = -32'd6264;
    weight_rom[102][34] = 32'd4802;
    weight_rom[102][35] = 32'd3694;
    weight_rom[102][36] = -32'd1062;
    weight_rom[102][37] = -32'd6031;
    weight_rom[102][38] = 32'd6124;
    weight_rom[102][39] = -32'd5961;
    weight_rom[102][40] = -32'd4351;
    weight_rom[102][41] = 32'd3056;
    weight_rom[102][42] = 32'd3489;
    weight_rom[102][43] = 32'd4845;
    weight_rom[102][44] = 32'd2321;
    weight_rom[102][45] = -32'd6455;
    weight_rom[102][46] = -32'd6379;
    weight_rom[102][47] = -32'd3079;
    weight_rom[102][48] = -32'd4367;
    weight_rom[102][49] = -32'd3809;
    weight_rom[102][50] = -32'd334;
    weight_rom[102][51] = -32'd1153;
    weight_rom[102][52] = 32'd6543;
    weight_rom[102][53] = -32'd3842;
    weight_rom[102][54] = 32'd55;
    weight_rom[102][55] = 32'd3600;
    weight_rom[102][56] = -32'd2349;
    weight_rom[102][57] = 32'd2438;
    weight_rom[102][58] = 32'd1119;
    weight_rom[102][59] = 32'd3308;
    weight_rom[102][60] = 32'd4970;
    weight_rom[102][61] = 32'd4989;
    weight_rom[102][62] = -32'd2012;
    weight_rom[102][63] = -32'd5868;
    weight_rom[103][0] = 32'd112;
    weight_rom[103][1] = 32'd34;
    weight_rom[103][2] = 32'd989;
    weight_rom[103][3] = -32'd2870;
    weight_rom[103][4] = 32'd5516;
    weight_rom[103][5] = 32'd35;
    weight_rom[103][6] = -32'd3004;
    weight_rom[103][7] = -32'd707;
    weight_rom[103][8] = -32'd1199;
    weight_rom[103][9] = -32'd913;
    weight_rom[103][10] = -32'd3170;
    weight_rom[103][11] = 32'd2859;
    weight_rom[103][12] = 32'd5596;
    weight_rom[103][13] = -32'd314;
    weight_rom[103][14] = 32'd3054;
    weight_rom[103][15] = -32'd5868;
    weight_rom[103][16] = -32'd4276;
    weight_rom[103][17] = -32'd5623;
    weight_rom[103][18] = -32'd3697;
    weight_rom[103][19] = 32'd4379;
    weight_rom[103][20] = 32'd2330;
    weight_rom[103][21] = 32'd6306;
    weight_rom[103][22] = -32'd2583;
    weight_rom[103][23] = -32'd2011;
    weight_rom[103][24] = -32'd4120;
    weight_rom[103][25] = -32'd2344;
    weight_rom[103][26] = 32'd6431;
    weight_rom[103][27] = -32'd529;
    weight_rom[103][28] = -32'd1476;
    weight_rom[103][29] = 32'd1017;
    weight_rom[103][30] = -32'd1401;
    weight_rom[103][31] = 32'd2313;
    weight_rom[103][32] = 32'd1534;
    weight_rom[103][33] = 32'd6324;
    weight_rom[103][34] = -32'd5772;
    weight_rom[103][35] = 32'd3484;
    weight_rom[103][36] = -32'd550;
    weight_rom[103][37] = -32'd2962;
    weight_rom[103][38] = 32'd2819;
    weight_rom[103][39] = -32'd813;
    weight_rom[103][40] = -32'd1903;
    weight_rom[103][41] = 32'd6493;
    weight_rom[103][42] = -32'd2567;
    weight_rom[103][43] = 32'd5122;
    weight_rom[103][44] = 32'd2394;
    weight_rom[103][45] = -32'd1013;
    weight_rom[103][46] = 32'd550;
    weight_rom[103][47] = 32'd2255;
    weight_rom[103][48] = 32'd3898;
    weight_rom[103][49] = -32'd6036;
    weight_rom[103][50] = -32'd6422;
    weight_rom[103][51] = -32'd4739;
    weight_rom[103][52] = -32'd2793;
    weight_rom[103][53] = -32'd1858;
    weight_rom[103][54] = 32'd4792;
    weight_rom[103][55] = -32'd3082;
    weight_rom[103][56] = 32'd6080;
    weight_rom[103][57] = -32'd3278;
    weight_rom[103][58] = 32'd624;
    weight_rom[103][59] = 32'd3320;
    weight_rom[103][60] = -32'd6383;
    weight_rom[103][61] = -32'd1141;
    weight_rom[103][62] = 32'd6200;
    weight_rom[103][63] = 32'd2431;
    weight_rom[104][0] = 32'd5342;
    weight_rom[104][1] = 32'd1008;
    weight_rom[104][2] = -32'd1465;
    weight_rom[104][3] = 32'd5903;
    weight_rom[104][4] = -32'd5753;
    weight_rom[104][5] = -32'd3509;
    weight_rom[104][6] = 32'd1887;
    weight_rom[104][7] = -32'd4126;
    weight_rom[104][8] = -32'd1668;
    weight_rom[104][9] = -32'd3925;
    weight_rom[104][10] = 32'd2054;
    weight_rom[104][11] = 32'd5970;
    weight_rom[104][12] = 32'd523;
    weight_rom[104][13] = -32'd1626;
    weight_rom[104][14] = 32'd1520;
    weight_rom[104][15] = -32'd1064;
    weight_rom[104][16] = 32'd2778;
    weight_rom[104][17] = -32'd3219;
    weight_rom[104][18] = 32'd6396;
    weight_rom[104][19] = 32'd3151;
    weight_rom[104][20] = 32'd1412;
    weight_rom[104][21] = 32'd911;
    weight_rom[104][22] = -32'd2289;
    weight_rom[104][23] = -32'd1342;
    weight_rom[104][24] = 32'd2152;
    weight_rom[104][25] = -32'd3668;
    weight_rom[104][26] = 32'd3365;
    weight_rom[104][27] = -32'd2536;
    weight_rom[104][28] = -32'd5686;
    weight_rom[104][29] = -32'd1845;
    weight_rom[104][30] = -32'd5239;
    weight_rom[104][31] = 32'd1235;
    weight_rom[104][32] = 32'd4586;
    weight_rom[104][33] = -32'd5424;
    weight_rom[104][34] = 32'd2517;
    weight_rom[104][35] = 32'd2512;
    weight_rom[104][36] = -32'd3189;
    weight_rom[104][37] = 32'd5972;
    weight_rom[104][38] = 32'd5991;
    weight_rom[104][39] = 32'd4508;
    weight_rom[104][40] = -32'd1310;
    weight_rom[104][41] = -32'd2785;
    weight_rom[104][42] = 32'd4084;
    weight_rom[104][43] = -32'd667;
    weight_rom[104][44] = 32'd1687;
    weight_rom[104][45] = 32'd2858;
    weight_rom[104][46] = -32'd529;
    weight_rom[104][47] = -32'd5871;
    weight_rom[104][48] = 32'd2885;
    weight_rom[104][49] = 32'd3162;
    weight_rom[104][50] = -32'd5442;
    weight_rom[104][51] = 32'd2172;
    weight_rom[104][52] = -32'd2877;
    weight_rom[104][53] = -32'd4595;
    weight_rom[104][54] = -32'd3390;
    weight_rom[104][55] = 32'd5683;
    weight_rom[104][56] = 32'd1855;
    weight_rom[104][57] = -32'd5693;
    weight_rom[104][58] = 32'd1841;
    weight_rom[104][59] = 32'd2835;
    weight_rom[104][60] = 32'd5829;
    weight_rom[104][61] = 32'd491;
    weight_rom[104][62] = 32'd6287;
    weight_rom[104][63] = -32'd836;
    weight_rom[105][0] = -32'd3286;
    weight_rom[105][1] = -32'd98;
    weight_rom[105][2] = 32'd1878;
    weight_rom[105][3] = 32'd5115;
    weight_rom[105][4] = -32'd2924;
    weight_rom[105][5] = 32'd5237;
    weight_rom[105][6] = -32'd1196;
    weight_rom[105][7] = 32'd549;
    weight_rom[105][8] = -32'd3148;
    weight_rom[105][9] = -32'd110;
    weight_rom[105][10] = -32'd2291;
    weight_rom[105][11] = -32'd6314;
    weight_rom[105][12] = 32'd4483;
    weight_rom[105][13] = -32'd1383;
    weight_rom[105][14] = -32'd4089;
    weight_rom[105][15] = -32'd3143;
    weight_rom[105][16] = 32'd4272;
    weight_rom[105][17] = -32'd1810;
    weight_rom[105][18] = -32'd602;
    weight_rom[105][19] = -32'd4681;
    weight_rom[105][20] = -32'd2683;
    weight_rom[105][21] = -32'd3151;
    weight_rom[105][22] = 32'd2786;
    weight_rom[105][23] = -32'd3089;
    weight_rom[105][24] = 32'd5002;
    weight_rom[105][25] = -32'd1959;
    weight_rom[105][26] = -32'd756;
    weight_rom[105][27] = 32'd4225;
    weight_rom[105][28] = -32'd6302;
    weight_rom[105][29] = 32'd4240;
    weight_rom[105][30] = -32'd6336;
    weight_rom[105][31] = 32'd1352;
    weight_rom[105][32] = -32'd3981;
    weight_rom[105][33] = 32'd4120;
    weight_rom[105][34] = -32'd4718;
    weight_rom[105][35] = 32'd6103;
    weight_rom[105][36] = 32'd3304;
    weight_rom[105][37] = 32'd5945;
    weight_rom[105][38] = -32'd955;
    weight_rom[105][39] = -32'd3114;
    weight_rom[105][40] = -32'd5801;
    weight_rom[105][41] = 32'd500;
    weight_rom[105][42] = -32'd2701;
    weight_rom[105][43] = -32'd533;
    weight_rom[105][44] = -32'd3065;
    weight_rom[105][45] = -32'd751;
    weight_rom[105][46] = -32'd13;
    weight_rom[105][47] = -32'd5064;
    weight_rom[105][48] = -32'd5424;
    weight_rom[105][49] = 32'd4294;
    weight_rom[105][50] = 32'd4032;
    weight_rom[105][51] = 32'd323;
    weight_rom[105][52] = -32'd4459;
    weight_rom[105][53] = 32'd130;
    weight_rom[105][54] = -32'd5524;
    weight_rom[105][55] = 32'd2883;
    weight_rom[105][56] = -32'd6246;
    weight_rom[105][57] = 32'd2498;
    weight_rom[105][58] = -32'd3152;
    weight_rom[105][59] = 32'd2220;
    weight_rom[105][60] = -32'd141;
    weight_rom[105][61] = -32'd5907;
    weight_rom[105][62] = -32'd3037;
    weight_rom[105][63] = -32'd4000;
    weight_rom[106][0] = -32'd1174;
    weight_rom[106][1] = -32'd3994;
    weight_rom[106][2] = -32'd547;
    weight_rom[106][3] = -32'd581;
    weight_rom[106][4] = 32'd4013;
    weight_rom[106][5] = -32'd1521;
    weight_rom[106][6] = -32'd6220;
    weight_rom[106][7] = 32'd4888;
    weight_rom[106][8] = 32'd2928;
    weight_rom[106][9] = -32'd5711;
    weight_rom[106][10] = 32'd3584;
    weight_rom[106][11] = -32'd3987;
    weight_rom[106][12] = 32'd274;
    weight_rom[106][13] = -32'd531;
    weight_rom[106][14] = -32'd1895;
    weight_rom[106][15] = 32'd3025;
    weight_rom[106][16] = -32'd5234;
    weight_rom[106][17] = -32'd360;
    weight_rom[106][18] = 32'd2467;
    weight_rom[106][19] = 32'd3321;
    weight_rom[106][20] = -32'd4763;
    weight_rom[106][21] = -32'd825;
    weight_rom[106][22] = 32'd4152;
    weight_rom[106][23] = -32'd3862;
    weight_rom[106][24] = 32'd4117;
    weight_rom[106][25] = -32'd1670;
    weight_rom[106][26] = 32'd2718;
    weight_rom[106][27] = -32'd5806;
    weight_rom[106][28] = 32'd4284;
    weight_rom[106][29] = 32'd4203;
    weight_rom[106][30] = 32'd2119;
    weight_rom[106][31] = 32'd2392;
    weight_rom[106][32] = -32'd4907;
    weight_rom[106][33] = -32'd2879;
    weight_rom[106][34] = -32'd1103;
    weight_rom[106][35] = -32'd1395;
    weight_rom[106][36] = 32'd168;
    weight_rom[106][37] = -32'd1935;
    weight_rom[106][38] = -32'd326;
    weight_rom[106][39] = -32'd1026;
    weight_rom[106][40] = 32'd1091;
    weight_rom[106][41] = 32'd436;
    weight_rom[106][42] = -32'd703;
    weight_rom[106][43] = -32'd5544;
    weight_rom[106][44] = -32'd6042;
    weight_rom[106][45] = 32'd3043;
    weight_rom[106][46] = -32'd5607;
    weight_rom[106][47] = -32'd6502;
    weight_rom[106][48] = -32'd474;
    weight_rom[106][49] = 32'd6132;
    weight_rom[106][50] = 32'd3558;
    weight_rom[106][51] = 32'd1826;
    weight_rom[106][52] = -32'd4403;
    weight_rom[106][53] = -32'd516;
    weight_rom[106][54] = -32'd1882;
    weight_rom[106][55] = 32'd3326;
    weight_rom[106][56] = -32'd915;
    weight_rom[106][57] = 32'd949;
    weight_rom[106][58] = -32'd5444;
    weight_rom[106][59] = -32'd301;
    weight_rom[106][60] = -32'd2071;
    weight_rom[106][61] = -32'd6522;
    weight_rom[106][62] = -32'd6016;
    weight_rom[106][63] = 32'd4142;
    weight_rom[107][0] = 32'd3349;
    weight_rom[107][1] = 32'd2915;
    weight_rom[107][2] = 32'd597;
    weight_rom[107][3] = 32'd1574;
    weight_rom[107][4] = 32'd3253;
    weight_rom[107][5] = 32'd570;
    weight_rom[107][6] = -32'd4506;
    weight_rom[107][7] = 32'd3043;
    weight_rom[107][8] = -32'd54;
    weight_rom[107][9] = 32'd1074;
    weight_rom[107][10] = -32'd4838;
    weight_rom[107][11] = -32'd6454;
    weight_rom[107][12] = 32'd1619;
    weight_rom[107][13] = 32'd3735;
    weight_rom[107][14] = 32'd3719;
    weight_rom[107][15] = 32'd6308;
    weight_rom[107][16] = -32'd3409;
    weight_rom[107][17] = -32'd5955;
    weight_rom[107][18] = -32'd4711;
    weight_rom[107][19] = 32'd3524;
    weight_rom[107][20] = 32'd1987;
    weight_rom[107][21] = 32'd1226;
    weight_rom[107][22] = -32'd4173;
    weight_rom[107][23] = -32'd222;
    weight_rom[107][24] = 32'd2426;
    weight_rom[107][25] = -32'd5652;
    weight_rom[107][26] = -32'd1451;
    weight_rom[107][27] = -32'd1066;
    weight_rom[107][28] = 32'd324;
    weight_rom[107][29] = -32'd296;
    weight_rom[107][30] = 32'd1342;
    weight_rom[107][31] = 32'd987;
    weight_rom[107][32] = 32'd6074;
    weight_rom[107][33] = -32'd4821;
    weight_rom[107][34] = 32'd636;
    weight_rom[107][35] = -32'd4840;
    weight_rom[107][36] = -32'd2348;
    weight_rom[107][37] = -32'd5988;
    weight_rom[107][38] = 32'd5216;
    weight_rom[107][39] = -32'd6030;
    weight_rom[107][40] = 32'd5037;
    weight_rom[107][41] = -32'd1236;
    weight_rom[107][42] = 32'd2975;
    weight_rom[107][43] = 32'd2238;
    weight_rom[107][44] = -32'd582;
    weight_rom[107][45] = -32'd3499;
    weight_rom[107][46] = 32'd2417;
    weight_rom[107][47] = 32'd6546;
    weight_rom[107][48] = -32'd4273;
    weight_rom[107][49] = 32'd5109;
    weight_rom[107][50] = 32'd5441;
    weight_rom[107][51] = -32'd2123;
    weight_rom[107][52] = -32'd2815;
    weight_rom[107][53] = 32'd5252;
    weight_rom[107][54] = 32'd3245;
    weight_rom[107][55] = -32'd3682;
    weight_rom[107][56] = 32'd4915;
    weight_rom[107][57] = -32'd1251;
    weight_rom[107][58] = -32'd4990;
    weight_rom[107][59] = 32'd1864;
    weight_rom[107][60] = 32'd5560;
    weight_rom[107][61] = -32'd3344;
    weight_rom[107][62] = 32'd2687;
    weight_rom[107][63] = 32'd3965;
    weight_rom[108][0] = -32'd3554;
    weight_rom[108][1] = -32'd2873;
    weight_rom[108][2] = 32'd5786;
    weight_rom[108][3] = -32'd2917;
    weight_rom[108][4] = -32'd4135;
    weight_rom[108][5] = 32'd5327;
    weight_rom[108][6] = 32'd2830;
    weight_rom[108][7] = 32'd4018;
    weight_rom[108][8] = -32'd5491;
    weight_rom[108][9] = -32'd3027;
    weight_rom[108][10] = 32'd6158;
    weight_rom[108][11] = 32'd1932;
    weight_rom[108][12] = -32'd5385;
    weight_rom[108][13] = 32'd5139;
    weight_rom[108][14] = 32'd710;
    weight_rom[108][15] = -32'd3191;
    weight_rom[108][16] = -32'd4692;
    weight_rom[108][17] = -32'd4718;
    weight_rom[108][18] = -32'd188;
    weight_rom[108][19] = 32'd2078;
    weight_rom[108][20] = 32'd3127;
    weight_rom[108][21] = -32'd5595;
    weight_rom[108][22] = -32'd1691;
    weight_rom[108][23] = -32'd3033;
    weight_rom[108][24] = -32'd5106;
    weight_rom[108][25] = -32'd1709;
    weight_rom[108][26] = -32'd3553;
    weight_rom[108][27] = -32'd544;
    weight_rom[108][28] = 32'd3607;
    weight_rom[108][29] = -32'd1955;
    weight_rom[108][30] = -32'd4416;
    weight_rom[108][31] = -32'd929;
    weight_rom[108][32] = -32'd5137;
    weight_rom[108][33] = -32'd788;
    weight_rom[108][34] = -32'd1274;
    weight_rom[108][35] = 32'd2250;
    weight_rom[108][36] = 32'd1258;
    weight_rom[108][37] = -32'd4206;
    weight_rom[108][38] = 32'd328;
    weight_rom[108][39] = -32'd667;
    weight_rom[108][40] = -32'd4564;
    weight_rom[108][41] = -32'd4336;
    weight_rom[108][42] = 32'd2528;
    weight_rom[108][43] = 32'd4210;
    weight_rom[108][44] = 32'd5124;
    weight_rom[108][45] = 32'd4104;
    weight_rom[108][46] = 32'd42;
    weight_rom[108][47] = 32'd3961;
    weight_rom[108][48] = -32'd2130;
    weight_rom[108][49] = 32'd1317;
    weight_rom[108][50] = 32'd4646;
    weight_rom[108][51] = 32'd5332;
    weight_rom[108][52] = 32'd3838;
    weight_rom[108][53] = 32'd5636;
    weight_rom[108][54] = 32'd664;
    weight_rom[108][55] = -32'd746;
    weight_rom[108][56] = -32'd2602;
    weight_rom[108][57] = -32'd1787;
    weight_rom[108][58] = -32'd3609;
    weight_rom[108][59] = -32'd6050;
    weight_rom[108][60] = -32'd6233;
    weight_rom[108][61] = 32'd2366;
    weight_rom[108][62] = -32'd642;
    weight_rom[108][63] = -32'd178;
    weight_rom[109][0] = -32'd5544;
    weight_rom[109][1] = -32'd6234;
    weight_rom[109][2] = -32'd1492;
    weight_rom[109][3] = -32'd4087;
    weight_rom[109][4] = -32'd3809;
    weight_rom[109][5] = 32'd1628;
    weight_rom[109][6] = 32'd2083;
    weight_rom[109][7] = 32'd2081;
    weight_rom[109][8] = -32'd3667;
    weight_rom[109][9] = 32'd3900;
    weight_rom[109][10] = -32'd605;
    weight_rom[109][11] = 32'd5217;
    weight_rom[109][12] = 32'd3345;
    weight_rom[109][13] = 32'd5968;
    weight_rom[109][14] = -32'd6485;
    weight_rom[109][15] = 32'd2020;
    weight_rom[109][16] = -32'd1993;
    weight_rom[109][17] = -32'd2925;
    weight_rom[109][18] = -32'd6192;
    weight_rom[109][19] = 32'd3488;
    weight_rom[109][20] = -32'd2416;
    weight_rom[109][21] = 32'd1603;
    weight_rom[109][22] = 32'd5268;
    weight_rom[109][23] = -32'd2785;
    weight_rom[109][24] = -32'd2763;
    weight_rom[109][25] = -32'd468;
    weight_rom[109][26] = 32'd1269;
    weight_rom[109][27] = 32'd2949;
    weight_rom[109][28] = -32'd3480;
    weight_rom[109][29] = -32'd1801;
    weight_rom[109][30] = -32'd3488;
    weight_rom[109][31] = -32'd2936;
    weight_rom[109][32] = -32'd281;
    weight_rom[109][33] = 32'd1886;
    weight_rom[109][34] = 32'd257;
    weight_rom[109][35] = 32'd3005;
    weight_rom[109][36] = 32'd6497;
    weight_rom[109][37] = -32'd1412;
    weight_rom[109][38] = 32'd2716;
    weight_rom[109][39] = 32'd1017;
    weight_rom[109][40] = 32'd1282;
    weight_rom[109][41] = 32'd6258;
    weight_rom[109][42] = 32'd6388;
    weight_rom[109][43] = -32'd3346;
    weight_rom[109][44] = 32'd910;
    weight_rom[109][45] = 32'd1159;
    weight_rom[109][46] = 32'd3475;
    weight_rom[109][47] = 32'd3758;
    weight_rom[109][48] = -32'd6316;
    weight_rom[109][49] = 32'd393;
    weight_rom[109][50] = 32'd2400;
    weight_rom[109][51] = 32'd1145;
    weight_rom[109][52] = 32'd5318;
    weight_rom[109][53] = -32'd1526;
    weight_rom[109][54] = 32'd4152;
    weight_rom[109][55] = 32'd1544;
    weight_rom[109][56] = -32'd5314;
    weight_rom[109][57] = -32'd3711;
    weight_rom[109][58] = 32'd2;
    weight_rom[109][59] = 32'd1592;
    weight_rom[109][60] = 32'd1067;
    weight_rom[109][61] = -32'd4964;
    weight_rom[109][62] = -32'd5232;
    weight_rom[109][63] = -32'd2641;
    weight_rom[110][0] = -32'd2755;
    weight_rom[110][1] = 32'd1906;
    weight_rom[110][2] = 32'd6044;
    weight_rom[110][3] = -32'd475;
    weight_rom[110][4] = -32'd1697;
    weight_rom[110][5] = -32'd5021;
    weight_rom[110][6] = -32'd6198;
    weight_rom[110][7] = 32'd2520;
    weight_rom[110][8] = 32'd2402;
    weight_rom[110][9] = -32'd2485;
    weight_rom[110][10] = -32'd3459;
    weight_rom[110][11] = -32'd3362;
    weight_rom[110][12] = -32'd4879;
    weight_rom[110][13] = 32'd3760;
    weight_rom[110][14] = 32'd3420;
    weight_rom[110][15] = -32'd3957;
    weight_rom[110][16] = -32'd650;
    weight_rom[110][17] = 32'd6180;
    weight_rom[110][18] = 32'd71;
    weight_rom[110][19] = 32'd4534;
    weight_rom[110][20] = 32'd1898;
    weight_rom[110][21] = 32'd6306;
    weight_rom[110][22] = 32'd4019;
    weight_rom[110][23] = 32'd2054;
    weight_rom[110][24] = -32'd2492;
    weight_rom[110][25] = 32'd2919;
    weight_rom[110][26] = 32'd5612;
    weight_rom[110][27] = 32'd973;
    weight_rom[110][28] = -32'd2030;
    weight_rom[110][29] = 32'd4007;
    weight_rom[110][30] = -32'd6242;
    weight_rom[110][31] = 32'd3520;
    weight_rom[110][32] = 32'd1121;
    weight_rom[110][33] = -32'd1560;
    weight_rom[110][34] = 32'd6508;
    weight_rom[110][35] = 32'd983;
    weight_rom[110][36] = -32'd848;
    weight_rom[110][37] = 32'd5869;
    weight_rom[110][38] = -32'd3248;
    weight_rom[110][39] = 32'd929;
    weight_rom[110][40] = 32'd2159;
    weight_rom[110][41] = 32'd4630;
    weight_rom[110][42] = -32'd3602;
    weight_rom[110][43] = -32'd1031;
    weight_rom[110][44] = 32'd4356;
    weight_rom[110][45] = -32'd3791;
    weight_rom[110][46] = -32'd192;
    weight_rom[110][47] = 32'd127;
    weight_rom[110][48] = -32'd1306;
    weight_rom[110][49] = -32'd6188;
    weight_rom[110][50] = -32'd5867;
    weight_rom[110][51] = -32'd5434;
    weight_rom[110][52] = 32'd6227;
    weight_rom[110][53] = -32'd108;
    weight_rom[110][54] = 32'd6023;
    weight_rom[110][55] = 32'd3538;
    weight_rom[110][56] = 32'd3386;
    weight_rom[110][57] = 32'd2223;
    weight_rom[110][58] = 32'd4462;
    weight_rom[110][59] = 32'd3642;
    weight_rom[110][60] = 32'd641;
    weight_rom[110][61] = -32'd5062;
    weight_rom[110][62] = 32'd2720;
    weight_rom[110][63] = 32'd1810;
    weight_rom[111][0] = -32'd4440;
    weight_rom[111][1] = -32'd4232;
    weight_rom[111][2] = 32'd5313;
    weight_rom[111][3] = -32'd1922;
    weight_rom[111][4] = -32'd202;
    weight_rom[111][5] = 32'd5764;
    weight_rom[111][6] = -32'd3644;
    weight_rom[111][7] = 32'd4576;
    weight_rom[111][8] = -32'd5555;
    weight_rom[111][9] = -32'd586;
    weight_rom[111][10] = -32'd5590;
    weight_rom[111][11] = 32'd5597;
    weight_rom[111][12] = 32'd4273;
    weight_rom[111][13] = -32'd2419;
    weight_rom[111][14] = -32'd6090;
    weight_rom[111][15] = 32'd856;
    weight_rom[111][16] = 32'd3261;
    weight_rom[111][17] = -32'd2210;
    weight_rom[111][18] = 32'd6081;
    weight_rom[111][19] = 32'd1489;
    weight_rom[111][20] = -32'd1374;
    weight_rom[111][21] = -32'd4061;
    weight_rom[111][22] = 32'd6355;
    weight_rom[111][23] = 32'd6141;
    weight_rom[111][24] = -32'd3277;
    weight_rom[111][25] = 32'd2054;
    weight_rom[111][26] = 32'd5624;
    weight_rom[111][27] = 32'd2191;
    weight_rom[111][28] = -32'd6159;
    weight_rom[111][29] = -32'd2252;
    weight_rom[111][30] = 32'd4390;
    weight_rom[111][31] = -32'd3587;
    weight_rom[111][32] = 32'd542;
    weight_rom[111][33] = -32'd5838;
    weight_rom[111][34] = -32'd4781;
    weight_rom[111][35] = -32'd3842;
    weight_rom[111][36] = 32'd5514;
    weight_rom[111][37] = -32'd4702;
    weight_rom[111][38] = -32'd698;
    weight_rom[111][39] = -32'd2196;
    weight_rom[111][40] = -32'd1057;
    weight_rom[111][41] = -32'd21;
    weight_rom[111][42] = 32'd2127;
    weight_rom[111][43] = 32'd4441;
    weight_rom[111][44] = 32'd6443;
    weight_rom[111][45] = -32'd3450;
    weight_rom[111][46] = -32'd4595;
    weight_rom[111][47] = -32'd2620;
    weight_rom[111][48] = 32'd653;
    weight_rom[111][49] = -32'd3320;
    weight_rom[111][50] = 32'd3707;
    weight_rom[111][51] = -32'd657;
    weight_rom[111][52] = -32'd3508;
    weight_rom[111][53] = 32'd5193;
    weight_rom[111][54] = 32'd3835;
    weight_rom[111][55] = -32'd5190;
    weight_rom[111][56] = 32'd1389;
    weight_rom[111][57] = 32'd6169;
    weight_rom[111][58] = 32'd2638;
    weight_rom[111][59] = 32'd4;
    weight_rom[111][60] = -32'd3678;
    weight_rom[111][61] = -32'd1167;
    weight_rom[111][62] = -32'd6144;
    weight_rom[111][63] = -32'd2776;
    weight_rom[112][0] = 32'd5632;
    weight_rom[112][1] = 32'd5773;
    weight_rom[112][2] = -32'd3987;
    weight_rom[112][3] = 32'd1096;
    weight_rom[112][4] = 32'd1549;
    weight_rom[112][5] = 32'd1673;
    weight_rom[112][6] = -32'd3524;
    weight_rom[112][7] = -32'd3281;
    weight_rom[112][8] = 32'd4603;
    weight_rom[112][9] = -32'd6401;
    weight_rom[112][10] = -32'd4328;
    weight_rom[112][11] = -32'd5763;
    weight_rom[112][12] = 32'd3696;
    weight_rom[112][13] = 32'd2465;
    weight_rom[112][14] = 32'd3220;
    weight_rom[112][15] = -32'd472;
    weight_rom[112][16] = 32'd1981;
    weight_rom[112][17] = -32'd235;
    weight_rom[112][18] = -32'd1517;
    weight_rom[112][19] = -32'd5392;
    weight_rom[112][20] = 32'd2794;
    weight_rom[112][21] = 32'd3835;
    weight_rom[112][22] = 32'd3332;
    weight_rom[112][23] = 32'd1358;
    weight_rom[112][24] = 32'd196;
    weight_rom[112][25] = 32'd2736;
    weight_rom[112][26] = -32'd2072;
    weight_rom[112][27] = 32'd3631;
    weight_rom[112][28] = 32'd6048;
    weight_rom[112][29] = -32'd3813;
    weight_rom[112][30] = 32'd6221;
    weight_rom[112][31] = 32'd2521;
    weight_rom[112][32] = -32'd5425;
    weight_rom[112][33] = 32'd1303;
    weight_rom[112][34] = 32'd2299;
    weight_rom[112][35] = 32'd58;
    weight_rom[112][36] = -32'd2031;
    weight_rom[112][37] = 32'd3453;
    weight_rom[112][38] = -32'd4935;
    weight_rom[112][39] = -32'd2417;
    weight_rom[112][40] = 32'd2635;
    weight_rom[112][41] = 32'd1353;
    weight_rom[112][42] = 32'd1437;
    weight_rom[112][43] = 32'd4942;
    weight_rom[112][44] = -32'd4409;
    weight_rom[112][45] = 32'd1678;
    weight_rom[112][46] = 32'd1943;
    weight_rom[112][47] = -32'd4570;
    weight_rom[112][48] = 32'd1567;
    weight_rom[112][49] = -32'd529;
    weight_rom[112][50] = 32'd4528;
    weight_rom[112][51] = 32'd3360;
    weight_rom[112][52] = 32'd4997;
    weight_rom[112][53] = 32'd4020;
    weight_rom[112][54] = 32'd1360;
    weight_rom[112][55] = 32'd6060;
    weight_rom[112][56] = 32'd921;
    weight_rom[112][57] = -32'd4250;
    weight_rom[112][58] = 32'd3788;
    weight_rom[112][59] = -32'd1867;
    weight_rom[112][60] = -32'd932;
    weight_rom[112][61] = 32'd1937;
    weight_rom[112][62] = 32'd4852;
    weight_rom[112][63] = -32'd3460;
    weight_rom[113][0] = 32'd4038;
    weight_rom[113][1] = 32'd5949;
    weight_rom[113][2] = -32'd5644;
    weight_rom[113][3] = -32'd5534;
    weight_rom[113][4] = -32'd1718;
    weight_rom[113][5] = -32'd2163;
    weight_rom[113][6] = 32'd2253;
    weight_rom[113][7] = -32'd138;
    weight_rom[113][8] = -32'd63;
    weight_rom[113][9] = -32'd5604;
    weight_rom[113][10] = 32'd259;
    weight_rom[113][11] = 32'd5694;
    weight_rom[113][12] = 32'd2736;
    weight_rom[113][13] = -32'd817;
    weight_rom[113][14] = -32'd3899;
    weight_rom[113][15] = 32'd6186;
    weight_rom[113][16] = 32'd1585;
    weight_rom[113][17] = -32'd3983;
    weight_rom[113][18] = -32'd6042;
    weight_rom[113][19] = -32'd162;
    weight_rom[113][20] = -32'd3942;
    weight_rom[113][21] = 32'd5346;
    weight_rom[113][22] = -32'd1399;
    weight_rom[113][23] = -32'd5544;
    weight_rom[113][24] = 32'd466;
    weight_rom[113][25] = -32'd6443;
    weight_rom[113][26] = 32'd362;
    weight_rom[113][27] = 32'd4747;
    weight_rom[113][28] = 32'd2200;
    weight_rom[113][29] = -32'd5443;
    weight_rom[113][30] = -32'd4778;
    weight_rom[113][31] = -32'd3495;
    weight_rom[113][32] = -32'd5806;
    weight_rom[113][33] = 32'd5274;
    weight_rom[113][34] = -32'd1363;
    weight_rom[113][35] = -32'd2461;
    weight_rom[113][36] = -32'd5836;
    weight_rom[113][37] = -32'd5129;
    weight_rom[113][38] = -32'd3853;
    weight_rom[113][39] = -32'd5156;
    weight_rom[113][40] = -32'd1170;
    weight_rom[113][41] = -32'd3574;
    weight_rom[113][42] = 32'd5440;
    weight_rom[113][43] = -32'd3366;
    weight_rom[113][44] = 32'd2513;
    weight_rom[113][45] = 32'd4324;
    weight_rom[113][46] = -32'd4294;
    weight_rom[113][47] = -32'd2822;
    weight_rom[113][48] = 32'd2142;
    weight_rom[113][49] = 32'd1684;
    weight_rom[113][50] = 32'd3920;
    weight_rom[113][51] = 32'd3855;
    weight_rom[113][52] = -32'd2251;
    weight_rom[113][53] = -32'd6505;
    weight_rom[113][54] = -32'd87;
    weight_rom[113][55] = 32'd5114;
    weight_rom[113][56] = -32'd5851;
    weight_rom[113][57] = 32'd1272;
    weight_rom[113][58] = -32'd1953;
    weight_rom[113][59] = -32'd2917;
    weight_rom[113][60] = 32'd1995;
    weight_rom[113][61] = 32'd2779;
    weight_rom[113][62] = -32'd4736;
    weight_rom[113][63] = 32'd3021;
    weight_rom[114][0] = 32'd1748;
    weight_rom[114][1] = 32'd5437;
    weight_rom[114][2] = -32'd5232;
    weight_rom[114][3] = 32'd6217;
    weight_rom[114][4] = -32'd491;
    weight_rom[114][5] = -32'd4728;
    weight_rom[114][6] = -32'd6295;
    weight_rom[114][7] = -32'd3654;
    weight_rom[114][8] = -32'd254;
    weight_rom[114][9] = -32'd1409;
    weight_rom[114][10] = -32'd2136;
    weight_rom[114][11] = -32'd1944;
    weight_rom[114][12] = -32'd6079;
    weight_rom[114][13] = -32'd3215;
    weight_rom[114][14] = 32'd6004;
    weight_rom[114][15] = 32'd1422;
    weight_rom[114][16] = -32'd1934;
    weight_rom[114][17] = 32'd1452;
    weight_rom[114][18] = -32'd6147;
    weight_rom[114][19] = -32'd5535;
    weight_rom[114][20] = 32'd5114;
    weight_rom[114][21] = 32'd5815;
    weight_rom[114][22] = 32'd1188;
    weight_rom[114][23] = -32'd5562;
    weight_rom[114][24] = -32'd1875;
    weight_rom[114][25] = -32'd3700;
    weight_rom[114][26] = -32'd3779;
    weight_rom[114][27] = -32'd2439;
    weight_rom[114][28] = 32'd5678;
    weight_rom[114][29] = -32'd436;
    weight_rom[114][30] = -32'd3519;
    weight_rom[114][31] = 32'd1642;
    weight_rom[114][32] = -32'd5170;
    weight_rom[114][33] = -32'd1530;
    weight_rom[114][34] = -32'd4810;
    weight_rom[114][35] = -32'd950;
    weight_rom[114][36] = -32'd3876;
    weight_rom[114][37] = 32'd6307;
    weight_rom[114][38] = -32'd6541;
    weight_rom[114][39] = -32'd1745;
    weight_rom[114][40] = 32'd60;
    weight_rom[114][41] = 32'd573;
    weight_rom[114][42] = -32'd4504;
    weight_rom[114][43] = 32'd662;
    weight_rom[114][44] = 32'd2284;
    weight_rom[114][45] = -32'd1105;
    weight_rom[114][46] = 32'd4881;
    weight_rom[114][47] = -32'd1625;
    weight_rom[114][48] = 32'd4407;
    weight_rom[114][49] = 32'd750;
    weight_rom[114][50] = 32'd111;
    weight_rom[114][51] = -32'd70;
    weight_rom[114][52] = -32'd5074;
    weight_rom[114][53] = -32'd2358;
    weight_rom[114][54] = -32'd6028;
    weight_rom[114][55] = -32'd3010;
    weight_rom[114][56] = -32'd4712;
    weight_rom[114][57] = -32'd993;
    weight_rom[114][58] = -32'd1249;
    weight_rom[114][59] = 32'd1871;
    weight_rom[114][60] = 32'd2977;
    weight_rom[114][61] = -32'd4214;
    weight_rom[114][62] = -32'd4884;
    weight_rom[114][63] = -32'd6025;
    weight_rom[115][0] = 32'd4868;
    weight_rom[115][1] = -32'd1701;
    weight_rom[115][2] = -32'd6314;
    weight_rom[115][3] = 32'd6372;
    weight_rom[115][4] = 32'd3243;
    weight_rom[115][5] = 32'd3853;
    weight_rom[115][6] = -32'd5189;
    weight_rom[115][7] = 32'd6391;
    weight_rom[115][8] = 32'd1211;
    weight_rom[115][9] = -32'd262;
    weight_rom[115][10] = 32'd4310;
    weight_rom[115][11] = -32'd5224;
    weight_rom[115][12] = -32'd2580;
    weight_rom[115][13] = 32'd4467;
    weight_rom[115][14] = -32'd1730;
    weight_rom[115][15] = -32'd1972;
    weight_rom[115][16] = 32'd4475;
    weight_rom[115][17] = -32'd2874;
    weight_rom[115][18] = -32'd1468;
    weight_rom[115][19] = -32'd1211;
    weight_rom[115][20] = -32'd2786;
    weight_rom[115][21] = 32'd6031;
    weight_rom[115][22] = 32'd2110;
    weight_rom[115][23] = 32'd5916;
    weight_rom[115][24] = -32'd1916;
    weight_rom[115][25] = 32'd2119;
    weight_rom[115][26] = 32'd6496;
    weight_rom[115][27] = 32'd498;
    weight_rom[115][28] = -32'd3073;
    weight_rom[115][29] = -32'd234;
    weight_rom[115][30] = 32'd4828;
    weight_rom[115][31] = 32'd3238;
    weight_rom[115][32] = 32'd1121;
    weight_rom[115][33] = -32'd3718;
    weight_rom[115][34] = -32'd4473;
    weight_rom[115][35] = 32'd1903;
    weight_rom[115][36] = -32'd1065;
    weight_rom[115][37] = -32'd1551;
    weight_rom[115][38] = -32'd6038;
    weight_rom[115][39] = -32'd5249;
    weight_rom[115][40] = -32'd6457;
    weight_rom[115][41] = 32'd2555;
    weight_rom[115][42] = 32'd3300;
    weight_rom[115][43] = -32'd4030;
    weight_rom[115][44] = 32'd6290;
    weight_rom[115][45] = -32'd3168;
    weight_rom[115][46] = 32'd1482;
    weight_rom[115][47] = 32'd3359;
    weight_rom[115][48] = -32'd3729;
    weight_rom[115][49] = 32'd3180;
    weight_rom[115][50] = -32'd3500;
    weight_rom[115][51] = 32'd5174;
    weight_rom[115][52] = 32'd4849;
    weight_rom[115][53] = -32'd1025;
    weight_rom[115][54] = 32'd6348;
    weight_rom[115][55] = 32'd4230;
    weight_rom[115][56] = 32'd1606;
    weight_rom[115][57] = -32'd698;
    weight_rom[115][58] = -32'd1393;
    weight_rom[115][59] = 32'd2527;
    weight_rom[115][60] = -32'd6544;
    weight_rom[115][61] = -32'd5510;
    weight_rom[115][62] = -32'd4251;
    weight_rom[115][63] = -32'd5311;
    weight_rom[116][0] = 32'd3980;
    weight_rom[116][1] = -32'd6351;
    weight_rom[116][2] = -32'd5315;
    weight_rom[116][3] = 32'd2597;
    weight_rom[116][4] = -32'd6072;
    weight_rom[116][5] = 32'd1573;
    weight_rom[116][6] = 32'd3931;
    weight_rom[116][7] = 32'd5820;
    weight_rom[116][8] = 32'd4255;
    weight_rom[116][9] = 32'd1310;
    weight_rom[116][10] = -32'd905;
    weight_rom[116][11] = -32'd185;
    weight_rom[116][12] = -32'd3104;
    weight_rom[116][13] = -32'd6049;
    weight_rom[116][14] = -32'd2268;
    weight_rom[116][15] = -32'd5058;
    weight_rom[116][16] = -32'd376;
    weight_rom[116][17] = -32'd3840;
    weight_rom[116][18] = -32'd4456;
    weight_rom[116][19] = -32'd1217;
    weight_rom[116][20] = -32'd1732;
    weight_rom[116][21] = 32'd281;
    weight_rom[116][22] = -32'd5525;
    weight_rom[116][23] = -32'd2656;
    weight_rom[116][24] = 32'd4306;
    weight_rom[116][25] = -32'd209;
    weight_rom[116][26] = 32'd6306;
    weight_rom[116][27] = 32'd4457;
    weight_rom[116][28] = 32'd1460;
    weight_rom[116][29] = 32'd4468;
    weight_rom[116][30] = 32'd5589;
    weight_rom[116][31] = -32'd3686;
    weight_rom[116][32] = 32'd581;
    weight_rom[116][33] = -32'd752;
    weight_rom[116][34] = 32'd5888;
    weight_rom[116][35] = 32'd3214;
    weight_rom[116][36] = -32'd3674;
    weight_rom[116][37] = 32'd3607;
    weight_rom[116][38] = 32'd6255;
    weight_rom[116][39] = 32'd3494;
    weight_rom[116][40] = 32'd2512;
    weight_rom[116][41] = 32'd198;
    weight_rom[116][42] = 32'd894;
    weight_rom[116][43] = -32'd5218;
    weight_rom[116][44] = 32'd6364;
    weight_rom[116][45] = 32'd4810;
    weight_rom[116][46] = -32'd4493;
    weight_rom[116][47] = 32'd519;
    weight_rom[116][48] = -32'd4974;
    weight_rom[116][49] = -32'd2886;
    weight_rom[116][50] = 32'd4526;
    weight_rom[116][51] = -32'd3045;
    weight_rom[116][52] = 32'd1783;
    weight_rom[116][53] = -32'd3542;
    weight_rom[116][54] = -32'd1527;
    weight_rom[116][55] = 32'd240;
    weight_rom[116][56] = -32'd3829;
    weight_rom[116][57] = -32'd3222;
    weight_rom[116][58] = -32'd4038;
    weight_rom[116][59] = 32'd4862;
    weight_rom[116][60] = 32'd5725;
    weight_rom[116][61] = 32'd5772;
    weight_rom[116][62] = 32'd6032;
    weight_rom[116][63] = -32'd6464;
    weight_rom[117][0] = -32'd4108;
    weight_rom[117][1] = 32'd5614;
    weight_rom[117][2] = 32'd2398;
    weight_rom[117][3] = 32'd473;
    weight_rom[117][4] = -32'd3244;
    weight_rom[117][5] = 32'd438;
    weight_rom[117][6] = -32'd4213;
    weight_rom[117][7] = -32'd6036;
    weight_rom[117][8] = -32'd1994;
    weight_rom[117][9] = -32'd2730;
    weight_rom[117][10] = -32'd3293;
    weight_rom[117][11] = -32'd3187;
    weight_rom[117][12] = -32'd1833;
    weight_rom[117][13] = 32'd5265;
    weight_rom[117][14] = -32'd4602;
    weight_rom[117][15] = -32'd4571;
    weight_rom[117][16] = 32'd6279;
    weight_rom[117][17] = 32'd217;
    weight_rom[117][18] = -32'd6247;
    weight_rom[117][19] = -32'd5688;
    weight_rom[117][20] = -32'd5792;
    weight_rom[117][21] = 32'd6256;
    weight_rom[117][22] = 32'd583;
    weight_rom[117][23] = -32'd5346;
    weight_rom[117][24] = 32'd3791;
    weight_rom[117][25] = -32'd6483;
    weight_rom[117][26] = 32'd1959;
    weight_rom[117][27] = 32'd6415;
    weight_rom[117][28] = 32'd2339;
    weight_rom[117][29] = -32'd3653;
    weight_rom[117][30] = -32'd1053;
    weight_rom[117][31] = -32'd5767;
    weight_rom[117][32] = -32'd3489;
    weight_rom[117][33] = -32'd5919;
    weight_rom[117][34] = 32'd4975;
    weight_rom[117][35] = -32'd3509;
    weight_rom[117][36] = -32'd6550;
    weight_rom[117][37] = -32'd2063;
    weight_rom[117][38] = -32'd3377;
    weight_rom[117][39] = 32'd6111;
    weight_rom[117][40] = 32'd2114;
    weight_rom[117][41] = 32'd6426;
    weight_rom[117][42] = -32'd2953;
    weight_rom[117][43] = 32'd5388;
    weight_rom[117][44] = 32'd2446;
    weight_rom[117][45] = 32'd2218;
    weight_rom[117][46] = 32'd6059;
    weight_rom[117][47] = -32'd5537;
    weight_rom[117][48] = 32'd4607;
    weight_rom[117][49] = 32'd851;
    weight_rom[117][50] = 32'd2977;
    weight_rom[117][51] = -32'd1171;
    weight_rom[117][52] = -32'd4394;
    weight_rom[117][53] = -32'd3937;
    weight_rom[117][54] = -32'd4558;
    weight_rom[117][55] = -32'd500;
    weight_rom[117][56] = 32'd53;
    weight_rom[117][57] = 32'd4261;
    weight_rom[117][58] = -32'd5751;
    weight_rom[117][59] = -32'd2066;
    weight_rom[117][60] = -32'd4397;
    weight_rom[117][61] = -32'd3137;
    weight_rom[117][62] = 32'd2531;
    weight_rom[117][63] = -32'd4548;
    weight_rom[118][0] = 32'd5145;
    weight_rom[118][1] = -32'd941;
    weight_rom[118][2] = -32'd5620;
    weight_rom[118][3] = -32'd2496;
    weight_rom[118][4] = 32'd2796;
    weight_rom[118][5] = 32'd5162;
    weight_rom[118][6] = 32'd2002;
    weight_rom[118][7] = 32'd2694;
    weight_rom[118][8] = 32'd2333;
    weight_rom[118][9] = 32'd2555;
    weight_rom[118][10] = 32'd1535;
    weight_rom[118][11] = -32'd2819;
    weight_rom[118][12] = -32'd5404;
    weight_rom[118][13] = -32'd504;
    weight_rom[118][14] = -32'd2547;
    weight_rom[118][15] = -32'd3600;
    weight_rom[118][16] = 32'd1758;
    weight_rom[118][17] = -32'd6481;
    weight_rom[118][18] = 32'd3358;
    weight_rom[118][19] = -32'd1981;
    weight_rom[118][20] = -32'd5092;
    weight_rom[118][21] = 32'd3372;
    weight_rom[118][22] = 32'd2743;
    weight_rom[118][23] = 32'd1298;
    weight_rom[118][24] = -32'd2519;
    weight_rom[118][25] = 32'd3991;
    weight_rom[118][26] = 32'd3990;
    weight_rom[118][27] = 32'd5105;
    weight_rom[118][28] = -32'd2391;
    weight_rom[118][29] = -32'd1559;
    weight_rom[118][30] = -32'd5890;
    weight_rom[118][31] = -32'd4836;
    weight_rom[118][32] = 32'd1805;
    weight_rom[118][33] = 32'd4200;
    weight_rom[118][34] = 32'd5335;
    weight_rom[118][35] = -32'd1240;
    weight_rom[118][36] = 32'd5439;
    weight_rom[118][37] = 32'd1673;
    weight_rom[118][38] = 32'd2140;
    weight_rom[118][39] = 32'd6161;
    weight_rom[118][40] = -32'd6050;
    weight_rom[118][41] = 32'd1459;
    weight_rom[118][42] = -32'd335;
    weight_rom[118][43] = 32'd4200;
    weight_rom[118][44] = -32'd3360;
    weight_rom[118][45] = -32'd680;
    weight_rom[118][46] = 32'd240;
    weight_rom[118][47] = -32'd6317;
    weight_rom[118][48] = -32'd4500;
    weight_rom[118][49] = -32'd5398;
    weight_rom[118][50] = 32'd6301;
    weight_rom[118][51] = 32'd5224;
    weight_rom[118][52] = -32'd919;
    weight_rom[118][53] = -32'd6058;
    weight_rom[118][54] = 32'd2185;
    weight_rom[118][55] = -32'd2432;
    weight_rom[118][56] = 32'd588;
    weight_rom[118][57] = -32'd193;
    weight_rom[118][58] = 32'd1191;
    weight_rom[118][59] = 32'd3535;
    weight_rom[118][60] = -32'd3492;
    weight_rom[118][61] = 32'd4631;
    weight_rom[118][62] = 32'd3950;
    weight_rom[118][63] = -32'd5649;
    weight_rom[119][0] = 32'd515;
    weight_rom[119][1] = 32'd6116;
    weight_rom[119][2] = -32'd2372;
    weight_rom[119][3] = 32'd4112;
    weight_rom[119][4] = 32'd5180;
    weight_rom[119][5] = 32'd3782;
    weight_rom[119][6] = -32'd3431;
    weight_rom[119][7] = 32'd5573;
    weight_rom[119][8] = 32'd861;
    weight_rom[119][9] = 32'd4720;
    weight_rom[119][10] = 32'd2710;
    weight_rom[119][11] = -32'd2525;
    weight_rom[119][12] = 32'd5727;
    weight_rom[119][13] = 32'd1798;
    weight_rom[119][14] = 32'd4936;
    weight_rom[119][15] = -32'd3264;
    weight_rom[119][16] = -32'd4898;
    weight_rom[119][17] = -32'd6453;
    weight_rom[119][18] = -32'd543;
    weight_rom[119][19] = -32'd5098;
    weight_rom[119][20] = 32'd207;
    weight_rom[119][21] = -32'd4434;
    weight_rom[119][22] = -32'd4360;
    weight_rom[119][23] = 32'd1620;
    weight_rom[119][24] = 32'd5423;
    weight_rom[119][25] = 32'd3575;
    weight_rom[119][26] = 32'd2819;
    weight_rom[119][27] = -32'd1684;
    weight_rom[119][28] = 32'd4562;
    weight_rom[119][29] = 32'd4042;
    weight_rom[119][30] = -32'd6037;
    weight_rom[119][31] = 32'd1389;
    weight_rom[119][32] = 32'd4195;
    weight_rom[119][33] = 32'd4277;
    weight_rom[119][34] = 32'd6442;
    weight_rom[119][35] = -32'd3025;
    weight_rom[119][36] = 32'd4507;
    weight_rom[119][37] = -32'd4036;
    weight_rom[119][38] = 32'd4444;
    weight_rom[119][39] = 32'd4785;
    weight_rom[119][40] = -32'd1726;
    weight_rom[119][41] = -32'd1691;
    weight_rom[119][42] = -32'd2178;
    weight_rom[119][43] = 32'd3408;
    weight_rom[119][44] = 32'd3913;
    weight_rom[119][45] = -32'd158;
    weight_rom[119][46] = -32'd5598;
    weight_rom[119][47] = -32'd5212;
    weight_rom[119][48] = 32'd6222;
    weight_rom[119][49] = -32'd1131;
    weight_rom[119][50] = -32'd4512;
    weight_rom[119][51] = 32'd5193;
    weight_rom[119][52] = -32'd2788;
    weight_rom[119][53] = 32'd1879;
    weight_rom[119][54] = -32'd2827;
    weight_rom[119][55] = 32'd1061;
    weight_rom[119][56] = -32'd2837;
    weight_rom[119][57] = 32'd568;
    weight_rom[119][58] = 32'd6412;
    weight_rom[119][59] = 32'd804;
    weight_rom[119][60] = -32'd3100;
    weight_rom[119][61] = 32'd4764;
    weight_rom[119][62] = -32'd1341;
    weight_rom[119][63] = 32'd6498;
    weight_rom[120][0] = 32'd4029;
    weight_rom[120][1] = 32'd6076;
    weight_rom[120][2] = 32'd4520;
    weight_rom[120][3] = 32'd2421;
    weight_rom[120][4] = 32'd153;
    weight_rom[120][5] = -32'd4565;
    weight_rom[120][6] = -32'd5250;
    weight_rom[120][7] = -32'd4186;
    weight_rom[120][8] = -32'd3053;
    weight_rom[120][9] = 32'd3668;
    weight_rom[120][10] = -32'd4364;
    weight_rom[120][11] = 32'd3971;
    weight_rom[120][12] = 32'd705;
    weight_rom[120][13] = 32'd2088;
    weight_rom[120][14] = 32'd6505;
    weight_rom[120][15] = 32'd4595;
    weight_rom[120][16] = 32'd2309;
    weight_rom[120][17] = -32'd3682;
    weight_rom[120][18] = -32'd2762;
    weight_rom[120][19] = 32'd4040;
    weight_rom[120][20] = -32'd3046;
    weight_rom[120][21] = -32'd302;
    weight_rom[120][22] = 32'd3678;
    weight_rom[120][23] = 32'd1946;
    weight_rom[120][24] = 32'd5935;
    weight_rom[120][25] = 32'd634;
    weight_rom[120][26] = 32'd1221;
    weight_rom[120][27] = -32'd3995;
    weight_rom[120][28] = 32'd5861;
    weight_rom[120][29] = 32'd4241;
    weight_rom[120][30] = 32'd969;
    weight_rom[120][31] = 32'd4580;
    weight_rom[120][32] = -32'd6008;
    weight_rom[120][33] = 32'd1153;
    weight_rom[120][34] = -32'd3823;
    weight_rom[120][35] = -32'd3950;
    weight_rom[120][36] = 32'd3175;
    weight_rom[120][37] = -32'd4639;
    weight_rom[120][38] = 32'd664;
    weight_rom[120][39] = 32'd1321;
    weight_rom[120][40] = 32'd6278;
    weight_rom[120][41] = 32'd3567;
    weight_rom[120][42] = 32'd1039;
    weight_rom[120][43] = -32'd5914;
    weight_rom[120][44] = -32'd5150;
    weight_rom[120][45] = -32'd3876;
    weight_rom[120][46] = 32'd1662;
    weight_rom[120][47] = -32'd1173;
    weight_rom[120][48] = 32'd4489;
    weight_rom[120][49] = 32'd3278;
    weight_rom[120][50] = -32'd3595;
    weight_rom[120][51] = 32'd2434;
    weight_rom[120][52] = 32'd3103;
    weight_rom[120][53] = -32'd3112;
    weight_rom[120][54] = 32'd1124;
    weight_rom[120][55] = 32'd3013;
    weight_rom[120][56] = 32'd5877;
    weight_rom[120][57] = -32'd2559;
    weight_rom[120][58] = -32'd4366;
    weight_rom[120][59] = 32'd5017;
    weight_rom[120][60] = -32'd6057;
    weight_rom[120][61] = 32'd3572;
    weight_rom[120][62] = -32'd2145;
    weight_rom[120][63] = -32'd2768;
    weight_rom[121][0] = 32'd5191;
    weight_rom[121][1] = 32'd4626;
    weight_rom[121][2] = -32'd6248;
    weight_rom[121][3] = -32'd4422;
    weight_rom[121][4] = 32'd420;
    weight_rom[121][5] = -32'd2467;
    weight_rom[121][6] = -32'd3366;
    weight_rom[121][7] = 32'd890;
    weight_rom[121][8] = 32'd4962;
    weight_rom[121][9] = -32'd6034;
    weight_rom[121][10] = -32'd4356;
    weight_rom[121][11] = 32'd513;
    weight_rom[121][12] = -32'd2549;
    weight_rom[121][13] = 32'd5178;
    weight_rom[121][14] = -32'd1726;
    weight_rom[121][15] = 32'd802;
    weight_rom[121][16] = -32'd2292;
    weight_rom[121][17] = -32'd6072;
    weight_rom[121][18] = 32'd5243;
    weight_rom[121][19] = 32'd5867;
    weight_rom[121][20] = 32'd4397;
    weight_rom[121][21] = 32'd2861;
    weight_rom[121][22] = 32'd1098;
    weight_rom[121][23] = -32'd3048;
    weight_rom[121][24] = -32'd2270;
    weight_rom[121][25] = -32'd5682;
    weight_rom[121][26] = -32'd5854;
    weight_rom[121][27] = -32'd139;
    weight_rom[121][28] = 32'd5044;
    weight_rom[121][29] = -32'd1512;
    weight_rom[121][30] = -32'd1403;
    weight_rom[121][31] = -32'd5963;
    weight_rom[121][32] = -32'd24;
    weight_rom[121][33] = -32'd1925;
    weight_rom[121][34] = -32'd1894;
    weight_rom[121][35] = 32'd3714;
    weight_rom[121][36] = -32'd4354;
    weight_rom[121][37] = 32'd5741;
    weight_rom[121][38] = -32'd4546;
    weight_rom[121][39] = 32'd2632;
    weight_rom[121][40] = -32'd1038;
    weight_rom[121][41] = -32'd4319;
    weight_rom[121][42] = 32'd5098;
    weight_rom[121][43] = 32'd4505;
    weight_rom[121][44] = 32'd3679;
    weight_rom[121][45] = 32'd1662;
    weight_rom[121][46] = -32'd3234;
    weight_rom[121][47] = 32'd5677;
    weight_rom[121][48] = 32'd11;
    weight_rom[121][49] = 32'd2534;
    weight_rom[121][50] = -32'd3777;
    weight_rom[121][51] = 32'd4705;
    weight_rom[121][52] = -32'd610;
    weight_rom[121][53] = -32'd5867;
    weight_rom[121][54] = 32'd1137;
    weight_rom[121][55] = -32'd1167;
    weight_rom[121][56] = 32'd4488;
    weight_rom[121][57] = -32'd4170;
    weight_rom[121][58] = -32'd5941;
    weight_rom[121][59] = 32'd364;
    weight_rom[121][60] = -32'd4940;
    weight_rom[121][61] = -32'd4340;
    weight_rom[121][62] = -32'd3480;
    weight_rom[121][63] = -32'd4597;
    weight_rom[122][0] = -32'd2385;
    weight_rom[122][1] = -32'd2694;
    weight_rom[122][2] = 32'd4121;
    weight_rom[122][3] = 32'd5386;
    weight_rom[122][4] = -32'd5148;
    weight_rom[122][5] = -32'd3296;
    weight_rom[122][6] = 32'd2913;
    weight_rom[122][7] = 32'd5445;
    weight_rom[122][8] = 32'd3898;
    weight_rom[122][9] = -32'd255;
    weight_rom[122][10] = -32'd6072;
    weight_rom[122][11] = -32'd2473;
    weight_rom[122][12] = -32'd1350;
    weight_rom[122][13] = 32'd1791;
    weight_rom[122][14] = -32'd673;
    weight_rom[122][15] = 32'd306;
    weight_rom[122][16] = 32'd2442;
    weight_rom[122][17] = -32'd5137;
    weight_rom[122][18] = -32'd5031;
    weight_rom[122][19] = -32'd5605;
    weight_rom[122][20] = -32'd6360;
    weight_rom[122][21] = -32'd3311;
    weight_rom[122][22] = 32'd5927;
    weight_rom[122][23] = -32'd6355;
    weight_rom[122][24] = -32'd1908;
    weight_rom[122][25] = 32'd3493;
    weight_rom[122][26] = -32'd592;
    weight_rom[122][27] = 32'd3167;
    weight_rom[122][28] = 32'd3133;
    weight_rom[122][29] = -32'd535;
    weight_rom[122][30] = -32'd6178;
    weight_rom[122][31] = 32'd3069;
    weight_rom[122][32] = 32'd2481;
    weight_rom[122][33] = 32'd3929;
    weight_rom[122][34] = 32'd2218;
    weight_rom[122][35] = 32'd5364;
    weight_rom[122][36] = -32'd4975;
    weight_rom[122][37] = 32'd5474;
    weight_rom[122][38] = 32'd2989;
    weight_rom[122][39] = -32'd2815;
    weight_rom[122][40] = 32'd25;
    weight_rom[122][41] = -32'd1513;
    weight_rom[122][42] = 32'd908;
    weight_rom[122][43] = -32'd812;
    weight_rom[122][44] = 32'd5376;
    weight_rom[122][45] = -32'd1851;
    weight_rom[122][46] = 32'd3980;
    weight_rom[122][47] = 32'd1800;
    weight_rom[122][48] = 32'd6310;
    weight_rom[122][49] = 32'd6430;
    weight_rom[122][50] = 32'd3834;
    weight_rom[122][51] = -32'd5390;
    weight_rom[122][52] = 32'd6413;
    weight_rom[122][53] = -32'd3526;
    weight_rom[122][54] = -32'd711;
    weight_rom[122][55] = 32'd1693;
    weight_rom[122][56] = 32'd2914;
    weight_rom[122][57] = -32'd5427;
    weight_rom[122][58] = 32'd3663;
    weight_rom[122][59] = 32'd231;
    weight_rom[122][60] = 32'd6374;
    weight_rom[122][61] = 32'd4217;
    weight_rom[122][62] = -32'd253;
    weight_rom[122][63] = -32'd3394;
    weight_rom[123][0] = -32'd5111;
    weight_rom[123][1] = -32'd1506;
    weight_rom[123][2] = -32'd2859;
    weight_rom[123][3] = 32'd4227;
    weight_rom[123][4] = -32'd689;
    weight_rom[123][5] = 32'd3197;
    weight_rom[123][6] = 32'd4662;
    weight_rom[123][7] = -32'd6108;
    weight_rom[123][8] = 32'd2076;
    weight_rom[123][9] = -32'd5178;
    weight_rom[123][10] = 32'd3098;
    weight_rom[123][11] = 32'd1446;
    weight_rom[123][12] = -32'd691;
    weight_rom[123][13] = 32'd1493;
    weight_rom[123][14] = 32'd2910;
    weight_rom[123][15] = -32'd5049;
    weight_rom[123][16] = -32'd5640;
    weight_rom[123][17] = -32'd2112;
    weight_rom[123][18] = 32'd5975;
    weight_rom[123][19] = 32'd5965;
    weight_rom[123][20] = -32'd1584;
    weight_rom[123][21] = 32'd1843;
    weight_rom[123][22] = -32'd5997;
    weight_rom[123][23] = 32'd6095;
    weight_rom[123][24] = 32'd73;
    weight_rom[123][25] = 32'd1097;
    weight_rom[123][26] = 32'd2290;
    weight_rom[123][27] = -32'd97;
    weight_rom[123][28] = -32'd2916;
    weight_rom[123][29] = -32'd2578;
    weight_rom[123][30] = 32'd1091;
    weight_rom[123][31] = -32'd2079;
    weight_rom[123][32] = -32'd3246;
    weight_rom[123][33] = 32'd716;
    weight_rom[123][34] = -32'd212;
    weight_rom[123][35] = -32'd1700;
    weight_rom[123][36] = -32'd5667;
    weight_rom[123][37] = 32'd5078;
    weight_rom[123][38] = 32'd1313;
    weight_rom[123][39] = 32'd1714;
    weight_rom[123][40] = 32'd5373;
    weight_rom[123][41] = -32'd2005;
    weight_rom[123][42] = 32'd1726;
    weight_rom[123][43] = -32'd2065;
    weight_rom[123][44] = -32'd1535;
    weight_rom[123][45] = 32'd6496;
    weight_rom[123][46] = 32'd4165;
    weight_rom[123][47] = 32'd3956;
    weight_rom[123][48] = -32'd5277;
    weight_rom[123][49] = -32'd2911;
    weight_rom[123][50] = -32'd4103;
    weight_rom[123][51] = 32'd4784;
    weight_rom[123][52] = -32'd5836;
    weight_rom[123][53] = 32'd3957;
    weight_rom[123][54] = 32'd4405;
    weight_rom[123][55] = 32'd2612;
    weight_rom[123][56] = -32'd5531;
    weight_rom[123][57] = 32'd2806;
    weight_rom[123][58] = -32'd3242;
    weight_rom[123][59] = 32'd1020;
    weight_rom[123][60] = -32'd2422;
    weight_rom[123][61] = 32'd3529;
    weight_rom[123][62] = 32'd679;
    weight_rom[123][63] = 32'd5716;
    weight_rom[124][0] = -32'd3566;
    weight_rom[124][1] = 32'd4602;
    weight_rom[124][2] = -32'd5004;
    weight_rom[124][3] = 32'd5895;
    weight_rom[124][4] = 32'd427;
    weight_rom[124][5] = -32'd6114;
    weight_rom[124][6] = 32'd4328;
    weight_rom[124][7] = 32'd2587;
    weight_rom[124][8] = 32'd4595;
    weight_rom[124][9] = -32'd3381;
    weight_rom[124][10] = 32'd2147;
    weight_rom[124][11] = 32'd2833;
    weight_rom[124][12] = 32'd1318;
    weight_rom[124][13] = -32'd5680;
    weight_rom[124][14] = 32'd5061;
    weight_rom[124][15] = 32'd4720;
    weight_rom[124][16] = -32'd4261;
    weight_rom[124][17] = 32'd3966;
    weight_rom[124][18] = -32'd2438;
    weight_rom[124][19] = 32'd295;
    weight_rom[124][20] = -32'd2131;
    weight_rom[124][21] = 32'd2183;
    weight_rom[124][22] = -32'd3075;
    weight_rom[124][23] = -32'd3265;
    weight_rom[124][24] = 32'd5781;
    weight_rom[124][25] = 32'd3695;
    weight_rom[124][26] = 32'd2326;
    weight_rom[124][27] = -32'd220;
    weight_rom[124][28] = -32'd2862;
    weight_rom[124][29] = 32'd5669;
    weight_rom[124][30] = -32'd6405;
    weight_rom[124][31] = -32'd281;
    weight_rom[124][32] = -32'd2519;
    weight_rom[124][33] = 32'd4272;
    weight_rom[124][34] = -32'd1069;
    weight_rom[124][35] = 32'd3293;
    weight_rom[124][36] = 32'd2936;
    weight_rom[124][37] = 32'd1644;
    weight_rom[124][38] = 32'd3031;
    weight_rom[124][39] = -32'd581;
    weight_rom[124][40] = 32'd2847;
    weight_rom[124][41] = -32'd893;
    weight_rom[124][42] = 32'd245;
    weight_rom[124][43] = 32'd609;
    weight_rom[124][44] = 32'd1712;
    weight_rom[124][45] = -32'd259;
    weight_rom[124][46] = 32'd6277;
    weight_rom[124][47] = -32'd440;
    weight_rom[124][48] = -32'd2581;
    weight_rom[124][49] = -32'd23;
    weight_rom[124][50] = -32'd5679;
    weight_rom[124][51] = -32'd2351;
    weight_rom[124][52] = -32'd1900;
    weight_rom[124][53] = 32'd4607;
    weight_rom[124][54] = -32'd3080;
    weight_rom[124][55] = 32'd2767;
    weight_rom[124][56] = -32'd5162;
    weight_rom[124][57] = -32'd3981;
    weight_rom[124][58] = 32'd4320;
    weight_rom[124][59] = 32'd3267;
    weight_rom[124][60] = -32'd5042;
    weight_rom[124][61] = 32'd1267;
    weight_rom[124][62] = 32'd1727;
    weight_rom[124][63] = 32'd264;
    weight_rom[125][0] = -32'd955;
    weight_rom[125][1] = -32'd2399;
    weight_rom[125][2] = 32'd2578;
    weight_rom[125][3] = 32'd2958;
    weight_rom[125][4] = -32'd3375;
    weight_rom[125][5] = 32'd916;
    weight_rom[125][6] = -32'd1347;
    weight_rom[125][7] = -32'd2656;
    weight_rom[125][8] = 32'd4814;
    weight_rom[125][9] = 32'd6378;
    weight_rom[125][10] = -32'd332;
    weight_rom[125][11] = -32'd2980;
    weight_rom[125][12] = 32'd205;
    weight_rom[125][13] = 32'd241;
    weight_rom[125][14] = 32'd1219;
    weight_rom[125][15] = 32'd2920;
    weight_rom[125][16] = 32'd4662;
    weight_rom[125][17] = 32'd944;
    weight_rom[125][18] = 32'd5090;
    weight_rom[125][19] = -32'd2627;
    weight_rom[125][20] = -32'd6300;
    weight_rom[125][21] = -32'd4421;
    weight_rom[125][22] = 32'd1331;
    weight_rom[125][23] = 32'd2307;
    weight_rom[125][24] = 32'd4932;
    weight_rom[125][25] = 32'd3299;
    weight_rom[125][26] = -32'd1662;
    weight_rom[125][27] = 32'd4433;
    weight_rom[125][28] = 32'd6073;
    weight_rom[125][29] = -32'd4998;
    weight_rom[125][30] = 32'd3766;
    weight_rom[125][31] = 32'd5621;
    weight_rom[125][32] = 32'd1489;
    weight_rom[125][33] = 32'd1723;
    weight_rom[125][34] = -32'd1863;
    weight_rom[125][35] = 32'd5203;
    weight_rom[125][36] = 32'd5620;
    weight_rom[125][37] = 32'd4040;
    weight_rom[125][38] = 32'd3535;
    weight_rom[125][39] = -32'd235;
    weight_rom[125][40] = 32'd1075;
    weight_rom[125][41] = 32'd3693;
    weight_rom[125][42] = -32'd5882;
    weight_rom[125][43] = -32'd5356;
    weight_rom[125][44] = -32'd915;
    weight_rom[125][45] = -32'd185;
    weight_rom[125][46] = 32'd24;
    weight_rom[125][47] = -32'd1813;
    weight_rom[125][48] = 32'd1811;
    weight_rom[125][49] = -32'd2234;
    weight_rom[125][50] = 32'd6534;
    weight_rom[125][51] = -32'd4216;
    weight_rom[125][52] = -32'd237;
    weight_rom[125][53] = -32'd221;
    weight_rom[125][54] = -32'd673;
    weight_rom[125][55] = -32'd5872;
    weight_rom[125][56] = -32'd94;
    weight_rom[125][57] = 32'd2491;
    weight_rom[125][58] = 32'd2673;
    weight_rom[125][59] = 32'd6090;
    weight_rom[125][60] = -32'd5151;
    weight_rom[125][61] = -32'd2133;
    weight_rom[125][62] = -32'd3183;
    weight_rom[125][63] = -32'd1771;
    weight_rom[126][0] = 32'd4168;
    weight_rom[126][1] = -32'd4331;
    weight_rom[126][2] = 32'd1690;
    weight_rom[126][3] = 32'd1486;
    weight_rom[126][4] = -32'd3024;
    weight_rom[126][5] = 32'd3440;
    weight_rom[126][6] = 32'd2203;
    weight_rom[126][7] = 32'd5562;
    weight_rom[126][8] = 32'd2731;
    weight_rom[126][9] = -32'd4685;
    weight_rom[126][10] = 32'd4511;
    weight_rom[126][11] = -32'd1133;
    weight_rom[126][12] = 32'd5497;
    weight_rom[126][13] = -32'd4585;
    weight_rom[126][14] = -32'd1421;
    weight_rom[126][15] = -32'd5666;
    weight_rom[126][16] = -32'd3575;
    weight_rom[126][17] = 32'd166;
    weight_rom[126][18] = 32'd1349;
    weight_rom[126][19] = -32'd5546;
    weight_rom[126][20] = -32'd4923;
    weight_rom[126][21] = 32'd853;
    weight_rom[126][22] = -32'd2666;
    weight_rom[126][23] = 32'd2708;
    weight_rom[126][24] = -32'd5209;
    weight_rom[126][25] = 32'd3971;
    weight_rom[126][26] = 32'd5789;
    weight_rom[126][27] = -32'd1816;
    weight_rom[126][28] = -32'd6418;
    weight_rom[126][29] = 32'd5685;
    weight_rom[126][30] = -32'd2537;
    weight_rom[126][31] = -32'd2202;
    weight_rom[126][32] = 32'd5215;
    weight_rom[126][33] = 32'd3727;
    weight_rom[126][34] = 32'd1229;
    weight_rom[126][35] = 32'd4536;
    weight_rom[126][36] = -32'd910;
    weight_rom[126][37] = -32'd5648;
    weight_rom[126][38] = 32'd6231;
    weight_rom[126][39] = 32'd3378;
    weight_rom[126][40] = 32'd3903;
    weight_rom[126][41] = -32'd207;
    weight_rom[126][42] = -32'd3501;
    weight_rom[126][43] = 32'd3363;
    weight_rom[126][44] = -32'd815;
    weight_rom[126][45] = 32'd863;
    weight_rom[126][46] = -32'd590;
    weight_rom[126][47] = -32'd5132;
    weight_rom[126][48] = -32'd1966;
    weight_rom[126][49] = -32'd778;
    weight_rom[126][50] = -32'd6228;
    weight_rom[126][51] = -32'd3416;
    weight_rom[126][52] = 32'd41;
    weight_rom[126][53] = -32'd1100;
    weight_rom[126][54] = 32'd494;
    weight_rom[126][55] = 32'd4715;
    weight_rom[126][56] = -32'd4447;
    weight_rom[126][57] = -32'd1436;
    weight_rom[126][58] = 32'd5841;
    weight_rom[126][59] = -32'd5589;
    weight_rom[126][60] = 32'd2876;
    weight_rom[126][61] = -32'd3112;
    weight_rom[126][62] = 32'd5880;
    weight_rom[126][63] = 32'd4894;
    weight_rom[127][0] = 32'd4728;
    weight_rom[127][1] = 32'd744;
    weight_rom[127][2] = 32'd4947;
    weight_rom[127][3] = -32'd1071;
    weight_rom[127][4] = -32'd1608;
    weight_rom[127][5] = 32'd4938;
    weight_rom[127][6] = -32'd3866;
    weight_rom[127][7] = 32'd6174;
    weight_rom[127][8] = 32'd4417;
    weight_rom[127][9] = -32'd14;
    weight_rom[127][10] = 32'd4006;
    weight_rom[127][11] = -32'd4956;
    weight_rom[127][12] = -32'd39;
    weight_rom[127][13] = 32'd3112;
    weight_rom[127][14] = -32'd1145;
    weight_rom[127][15] = 32'd2724;
    weight_rom[127][16] = 32'd4417;
    weight_rom[127][17] = -32'd2706;
    weight_rom[127][18] = 32'd4282;
    weight_rom[127][19] = 32'd8;
    weight_rom[127][20] = -32'd1131;
    weight_rom[127][21] = 32'd3560;
    weight_rom[127][22] = 32'd2810;
    weight_rom[127][23] = 32'd1441;
    weight_rom[127][24] = -32'd1406;
    weight_rom[127][25] = 32'd236;
    weight_rom[127][26] = -32'd4360;
    weight_rom[127][27] = 32'd4715;
    weight_rom[127][28] = 32'd2831;
    weight_rom[127][29] = 32'd2409;
    weight_rom[127][30] = -32'd6025;
    weight_rom[127][31] = -32'd454;
    weight_rom[127][32] = 32'd4062;
    weight_rom[127][33] = 32'd1291;
    weight_rom[127][34] = 32'd990;
    weight_rom[127][35] = -32'd4157;
    weight_rom[127][36] = -32'd4992;
    weight_rom[127][37] = -32'd2165;
    weight_rom[127][38] = 32'd964;
    weight_rom[127][39] = -32'd2858;
    weight_rom[127][40] = 32'd4775;
    weight_rom[127][41] = 32'd3853;
    weight_rom[127][42] = -32'd104;
    weight_rom[127][43] = 32'd1080;
    weight_rom[127][44] = -32'd2485;
    weight_rom[127][45] = 32'd5462;
    weight_rom[127][46] = 32'd3322;
    weight_rom[127][47] = 32'd4927;
    weight_rom[127][48] = 32'd5614;
    weight_rom[127][49] = 32'd4678;
    weight_rom[127][50] = 32'd4394;
    weight_rom[127][51] = -32'd1075;
    weight_rom[127][52] = -32'd2412;
    weight_rom[127][53] = 32'd6263;
    weight_rom[127][54] = 32'd2144;
    weight_rom[127][55] = -32'd547;
    weight_rom[127][56] = 32'd6268;
    weight_rom[127][57] = -32'd1103;
    weight_rom[127][58] = -32'd1193;
    weight_rom[127][59] = -32'd5853;
    weight_rom[127][60] = 32'd4647;
    weight_rom[127][61] = -32'd4955;
    weight_rom[127][62] = -32'd4328;
    weight_rom[127][63] = -32'd1376;
//end
// Initialization of biases
//initial begin
    bias_rom[0] = -32'd2162;
    bias_rom[1] = -32'd3836;
    bias_rom[2] = -32'd1601;
    bias_rom[3] = -32'd2402;
    bias_rom[4] = 32'd2323;
    bias_rom[5] = -32'd2757;
    bias_rom[6] = 32'd1011;
    bias_rom[7] = -32'd5689;
    bias_rom[8] = -32'd4046;
    bias_rom[9] = -32'd1213;
    bias_rom[10] = 32'd5727;
    bias_rom[11] = -32'd1608;
    bias_rom[12] = 32'd2150;
    bias_rom[13] = -32'd3210;
    bias_rom[14] = -32'd4888;
    bias_rom[15] = -32'd5786;
    bias_rom[16] = -32'd2550;
    bias_rom[17] = -32'd4487;
    bias_rom[18] = -32'd4272;
    bias_rom[19] = 32'd3417;
    bias_rom[20] = -32'd6345;
    bias_rom[21] = 32'd757;
    bias_rom[22] = -32'd1579;
    bias_rom[23] = 32'd85;
    bias_rom[24] = 32'd823;
    bias_rom[25] = -32'd2446;
    bias_rom[26] = -32'd2685;
    bias_rom[27] = 32'd3059;
    bias_rom[28] = 32'd4866;
    bias_rom[29] = -32'd4029;
    bias_rom[30] = -32'd5274;
    bias_rom[31] = 32'd5213;
    bias_rom[32] = -32'd1967;
    bias_rom[33] = 32'd672;
    bias_rom[34] = -32'd1840;
    bias_rom[35] = -32'd4904;
    bias_rom[36] = 32'd1170;
    bias_rom[37] = 32'd329;
    bias_rom[38] = -32'd3892;
    bias_rom[39] = -32'd630;
    bias_rom[40] = 32'd3892;
    bias_rom[41] = 32'd1185;
    bias_rom[42] = -32'd5283;
    bias_rom[43] = 32'd629;
    bias_rom[44] = 32'd2657;
    bias_rom[45] = 32'd3836;
    bias_rom[46] = 32'd1692;
    bias_rom[47] = -32'd4552;
    bias_rom[48] = 32'd2754;
    bias_rom[49] = 32'd2324;
    bias_rom[50] = -32'd6233;
    bias_rom[51] = -32'd1156;
    bias_rom[52] = -32'd2189;
    bias_rom[53] = 32'd2220;
    bias_rom[54] = -32'd3720;
    bias_rom[55] = 32'd1191;
    bias_rom[56] = 32'd5415;
    bias_rom[57] = 32'd3903;
    bias_rom[58] = 32'd5524;
    bias_rom[59] = 32'd6271;
    bias_rom[60] = -32'd6413;
    bias_rom[61] = 32'd1608;
    bias_rom[62] = -32'd1142;
    bias_rom[63] = 32'd4716;
//end
endtask
